
module CacheController ( rst, clk, wr, rd, data_rd, data_wr, addr_req, 
        addr_resp, rdy, busy, wr_mem, rd_mem, busy_mem, data_rd_mem, 
        data_wr_mem, addr_mem, cache_miss_count, cache_hit_count );
  output [31:0] data_rd;
  input [31:0] data_wr;
  input [31:0] addr_req;
  output [31:0] addr_resp;
  input [31:0] data_rd_mem;
  output [31:0] data_wr_mem;
  output [31:0] addr_mem;
  output [31:0] cache_miss_count;
  output [31:0] cache_hit_count;
  input rst, clk, wr, rd, busy_mem;
  output rdy, busy, wr_mem, rd_mem;
  wire   valid, dirty, miss, mem_done, hit, \cache_tag[15][23] ,
         \cache_tag[15][22] , \cache_tag[15][21] , \cache_tag[15][20] ,
         \cache_tag[15][19] , \cache_tag[15][18] , \cache_tag[15][17] ,
         \cache_tag[15][16] , \cache_tag[15][15] , \cache_tag[15][14] ,
         \cache_tag[15][13] , \cache_tag[15][12] , \cache_tag[15][11] ,
         \cache_tag[15][10] , \cache_tag[15][9] , \cache_tag[15][8] ,
         \cache_tag[15][7] , \cache_tag[15][6] , \cache_tag[15][5] ,
         \cache_tag[15][4] , \cache_tag[15][3] , \cache_tag[15][2] ,
         \cache_tag[15][1] , \cache_tag[15][0] , \cache_tag[14][23] ,
         \cache_tag[14][22] , \cache_tag[14][21] , \cache_tag[14][20] ,
         \cache_tag[14][19] , \cache_tag[14][18] , \cache_tag[14][17] ,
         \cache_tag[14][16] , \cache_tag[14][15] , \cache_tag[14][14] ,
         \cache_tag[14][13] , \cache_tag[14][12] , \cache_tag[14][11] ,
         \cache_tag[14][10] , \cache_tag[14][9] , \cache_tag[14][8] ,
         \cache_tag[14][7] , \cache_tag[14][6] , \cache_tag[14][5] ,
         \cache_tag[14][4] , \cache_tag[14][3] , \cache_tag[14][2] ,
         \cache_tag[14][1] , \cache_tag[14][0] , \cache_tag[13][23] ,
         \cache_tag[13][22] , \cache_tag[13][21] , \cache_tag[13][20] ,
         \cache_tag[13][19] , \cache_tag[13][18] , \cache_tag[13][17] ,
         \cache_tag[13][16] , \cache_tag[13][15] , \cache_tag[13][14] ,
         \cache_tag[13][13] , \cache_tag[13][12] , \cache_tag[13][11] ,
         \cache_tag[13][10] , \cache_tag[13][9] , \cache_tag[13][8] ,
         \cache_tag[13][7] , \cache_tag[13][6] , \cache_tag[13][5] ,
         \cache_tag[13][4] , \cache_tag[13][3] , \cache_tag[13][2] ,
         \cache_tag[13][1] , \cache_tag[13][0] , \cache_tag[12][23] ,
         \cache_tag[12][22] , \cache_tag[12][21] , \cache_tag[12][20] ,
         \cache_tag[12][19] , \cache_tag[12][18] , \cache_tag[12][17] ,
         \cache_tag[12][16] , \cache_tag[12][15] , \cache_tag[12][14] ,
         \cache_tag[12][13] , \cache_tag[12][12] , \cache_tag[12][11] ,
         \cache_tag[12][10] , \cache_tag[12][9] , \cache_tag[12][8] ,
         \cache_tag[12][7] , \cache_tag[12][6] , \cache_tag[12][5] ,
         \cache_tag[12][4] , \cache_tag[12][3] , \cache_tag[12][2] ,
         \cache_tag[12][1] , \cache_tag[12][0] , \cache_tag[11][23] ,
         \cache_tag[11][22] , \cache_tag[11][21] , \cache_tag[11][20] ,
         \cache_tag[11][19] , \cache_tag[11][18] , \cache_tag[11][17] ,
         \cache_tag[11][16] , \cache_tag[11][15] , \cache_tag[11][14] ,
         \cache_tag[11][13] , \cache_tag[11][12] , \cache_tag[11][11] ,
         \cache_tag[11][10] , \cache_tag[11][9] , \cache_tag[11][8] ,
         \cache_tag[11][7] , \cache_tag[11][6] , \cache_tag[11][5] ,
         \cache_tag[11][4] , \cache_tag[11][3] , \cache_tag[11][2] ,
         \cache_tag[11][1] , \cache_tag[11][0] , \cache_tag[10][23] ,
         \cache_tag[10][22] , \cache_tag[10][21] , \cache_tag[10][20] ,
         \cache_tag[10][19] , \cache_tag[10][18] , \cache_tag[10][17] ,
         \cache_tag[10][16] , \cache_tag[10][15] , \cache_tag[10][14] ,
         \cache_tag[10][13] , \cache_tag[10][12] , \cache_tag[10][11] ,
         \cache_tag[10][10] , \cache_tag[10][9] , \cache_tag[10][8] ,
         \cache_tag[10][7] , \cache_tag[10][6] , \cache_tag[10][5] ,
         \cache_tag[10][4] , \cache_tag[10][3] , \cache_tag[10][2] ,
         \cache_tag[10][1] , \cache_tag[10][0] , \cache_tag[9][23] ,
         \cache_tag[9][22] , \cache_tag[9][21] , \cache_tag[9][20] ,
         \cache_tag[9][19] , \cache_tag[9][18] , \cache_tag[9][17] ,
         \cache_tag[9][16] , \cache_tag[9][15] , \cache_tag[9][14] ,
         \cache_tag[9][13] , \cache_tag[9][12] , \cache_tag[9][11] ,
         \cache_tag[9][10] , \cache_tag[9][9] , \cache_tag[9][8] ,
         \cache_tag[9][7] , \cache_tag[9][6] , \cache_tag[9][5] ,
         \cache_tag[9][4] , \cache_tag[9][3] , \cache_tag[9][2] ,
         \cache_tag[9][1] , \cache_tag[9][0] , \cache_tag[8][23] ,
         \cache_tag[8][22] , \cache_tag[8][21] , \cache_tag[8][20] ,
         \cache_tag[8][19] , \cache_tag[8][18] , \cache_tag[8][17] ,
         \cache_tag[8][16] , \cache_tag[8][15] , \cache_tag[8][14] ,
         \cache_tag[8][13] , \cache_tag[8][12] , \cache_tag[8][11] ,
         \cache_tag[8][10] , \cache_tag[8][9] , \cache_tag[8][8] ,
         \cache_tag[8][7] , \cache_tag[8][6] , \cache_tag[8][5] ,
         \cache_tag[8][4] , \cache_tag[8][3] , \cache_tag[8][2] ,
         \cache_tag[8][1] , \cache_tag[8][0] , \cache_tag[7][23] ,
         \cache_tag[7][22] , \cache_tag[7][21] , \cache_tag[7][20] ,
         \cache_tag[7][19] , \cache_tag[7][18] , \cache_tag[7][17] ,
         \cache_tag[7][16] , \cache_tag[7][15] , \cache_tag[7][14] ,
         \cache_tag[7][13] , \cache_tag[7][12] , \cache_tag[7][11] ,
         \cache_tag[7][10] , \cache_tag[7][9] , \cache_tag[7][8] ,
         \cache_tag[7][7] , \cache_tag[7][6] , \cache_tag[7][5] ,
         \cache_tag[7][4] , \cache_tag[7][3] , \cache_tag[7][2] ,
         \cache_tag[7][1] , \cache_tag[7][0] , \cache_tag[6][23] ,
         \cache_tag[6][22] , \cache_tag[6][21] , \cache_tag[6][20] ,
         \cache_tag[6][19] , \cache_tag[6][18] , \cache_tag[6][17] ,
         \cache_tag[6][16] , \cache_tag[6][15] , \cache_tag[6][14] ,
         \cache_tag[6][13] , \cache_tag[6][12] , \cache_tag[6][11] ,
         \cache_tag[6][10] , \cache_tag[6][9] , \cache_tag[6][8] ,
         \cache_tag[6][7] , \cache_tag[6][6] , \cache_tag[6][5] ,
         \cache_tag[6][4] , \cache_tag[6][3] , \cache_tag[6][2] ,
         \cache_tag[6][1] , \cache_tag[6][0] , \cache_tag[5][23] ,
         \cache_tag[5][22] , \cache_tag[5][21] , \cache_tag[5][20] ,
         \cache_tag[5][19] , \cache_tag[5][18] , \cache_tag[5][17] ,
         \cache_tag[5][16] , \cache_tag[5][15] , \cache_tag[5][14] ,
         \cache_tag[5][13] , \cache_tag[5][12] , \cache_tag[5][11] ,
         \cache_tag[5][10] , \cache_tag[5][9] , \cache_tag[5][8] ,
         \cache_tag[5][7] , \cache_tag[5][6] , \cache_tag[5][5] ,
         \cache_tag[5][4] , \cache_tag[5][3] , \cache_tag[5][2] ,
         \cache_tag[5][1] , \cache_tag[5][0] , \cache_tag[4][23] ,
         \cache_tag[4][22] , \cache_tag[4][21] , \cache_tag[4][20] ,
         \cache_tag[4][19] , \cache_tag[4][18] , \cache_tag[4][17] ,
         \cache_tag[4][16] , \cache_tag[4][15] , \cache_tag[4][14] ,
         \cache_tag[4][13] , \cache_tag[4][12] , \cache_tag[4][11] ,
         \cache_tag[4][10] , \cache_tag[4][9] , \cache_tag[4][8] ,
         \cache_tag[4][7] , \cache_tag[4][6] , \cache_tag[4][5] ,
         \cache_tag[4][4] , \cache_tag[4][3] , \cache_tag[4][2] ,
         \cache_tag[4][1] , \cache_tag[4][0] , \cache_tag[3][23] ,
         \cache_tag[3][22] , \cache_tag[3][21] , \cache_tag[3][20] ,
         \cache_tag[3][19] , \cache_tag[3][18] , \cache_tag[3][17] ,
         \cache_tag[3][16] , \cache_tag[3][15] , \cache_tag[3][14] ,
         \cache_tag[3][13] , \cache_tag[3][12] , \cache_tag[3][11] ,
         \cache_tag[3][10] , \cache_tag[3][9] , \cache_tag[3][8] ,
         \cache_tag[3][7] , \cache_tag[3][6] , \cache_tag[3][5] ,
         \cache_tag[3][4] , \cache_tag[3][3] , \cache_tag[3][2] ,
         \cache_tag[3][1] , \cache_tag[3][0] , \cache_tag[2][23] ,
         \cache_tag[2][22] , \cache_tag[2][21] , \cache_tag[2][20] ,
         \cache_tag[2][19] , \cache_tag[2][18] , \cache_tag[2][17] ,
         \cache_tag[2][16] , \cache_tag[2][15] , \cache_tag[2][14] ,
         \cache_tag[2][13] , \cache_tag[2][12] , \cache_tag[2][11] ,
         \cache_tag[2][10] , \cache_tag[2][9] , \cache_tag[2][8] ,
         \cache_tag[2][7] , \cache_tag[2][6] , \cache_tag[2][5] ,
         \cache_tag[2][4] , \cache_tag[2][3] , \cache_tag[2][2] ,
         \cache_tag[2][1] , \cache_tag[2][0] , \cache_tag[1][23] ,
         \cache_tag[1][22] , \cache_tag[1][21] , \cache_tag[1][20] ,
         \cache_tag[1][19] , \cache_tag[1][18] , \cache_tag[1][17] ,
         \cache_tag[1][16] , \cache_tag[1][15] , \cache_tag[1][14] ,
         \cache_tag[1][13] , \cache_tag[1][12] , \cache_tag[1][11] ,
         \cache_tag[1][10] , \cache_tag[1][9] , \cache_tag[1][8] ,
         \cache_tag[1][7] , \cache_tag[1][6] , \cache_tag[1][5] ,
         \cache_tag[1][4] , \cache_tag[1][3] , \cache_tag[1][2] ,
         \cache_tag[1][1] , \cache_tag[1][0] , \cache_tag[0][23] ,
         \cache_tag[0][22] , \cache_tag[0][21] , \cache_tag[0][20] ,
         \cache_tag[0][19] , \cache_tag[0][18] , \cache_tag[0][17] ,
         \cache_tag[0][16] , \cache_tag[0][15] , \cache_tag[0][14] ,
         \cache_tag[0][13] , \cache_tag[0][12] , \cache_tag[0][11] ,
         \cache_tag[0][10] , \cache_tag[0][9] , \cache_tag[0][8] ,
         \cache_tag[0][7] , \cache_tag[0][6] , \cache_tag[0][5] ,
         \cache_tag[0][4] , \cache_tag[0][3] , \cache_tag[0][2] ,
         \cache_tag[0][1] , \cache_tag[0][0] , \cache_data[15][127] ,
         \cache_data[15][126] , \cache_data[15][125] , \cache_data[15][124] ,
         \cache_data[15][123] , \cache_data[15][122] , \cache_data[15][121] ,
         \cache_data[15][120] , \cache_data[15][119] , \cache_data[15][118] ,
         \cache_data[15][117] , \cache_data[15][116] , \cache_data[15][115] ,
         \cache_data[15][114] , \cache_data[15][113] , \cache_data[15][112] ,
         \cache_data[15][111] , \cache_data[15][110] , \cache_data[15][109] ,
         \cache_data[15][108] , \cache_data[15][107] , \cache_data[15][106] ,
         \cache_data[15][105] , \cache_data[15][104] , \cache_data[15][103] ,
         \cache_data[15][102] , \cache_data[15][101] , \cache_data[15][100] ,
         \cache_data[15][99] , \cache_data[15][98] , \cache_data[15][97] ,
         \cache_data[15][96] , \cache_data[15][95] , \cache_data[15][94] ,
         \cache_data[15][93] , \cache_data[15][92] , \cache_data[15][91] ,
         \cache_data[15][90] , \cache_data[15][89] , \cache_data[15][88] ,
         \cache_data[15][87] , \cache_data[15][86] , \cache_data[15][85] ,
         \cache_data[15][84] , \cache_data[15][83] , \cache_data[15][82] ,
         \cache_data[15][81] , \cache_data[15][80] , \cache_data[15][79] ,
         \cache_data[15][78] , \cache_data[15][77] , \cache_data[15][76] ,
         \cache_data[15][75] , \cache_data[15][74] , \cache_data[15][73] ,
         \cache_data[15][72] , \cache_data[15][71] , \cache_data[15][70] ,
         \cache_data[15][69] , \cache_data[15][68] , \cache_data[15][67] ,
         \cache_data[15][66] , \cache_data[15][65] , \cache_data[15][64] ,
         \cache_data[15][63] , \cache_data[15][62] , \cache_data[15][61] ,
         \cache_data[15][60] , \cache_data[15][59] , \cache_data[15][58] ,
         \cache_data[15][57] , \cache_data[15][56] , \cache_data[15][55] ,
         \cache_data[15][54] , \cache_data[15][53] , \cache_data[15][52] ,
         \cache_data[15][51] , \cache_data[15][50] , \cache_data[15][49] ,
         \cache_data[15][48] , \cache_data[15][47] , \cache_data[15][46] ,
         \cache_data[15][45] , \cache_data[15][44] , \cache_data[15][43] ,
         \cache_data[15][42] , \cache_data[15][41] , \cache_data[15][40] ,
         \cache_data[15][39] , \cache_data[15][38] , \cache_data[15][37] ,
         \cache_data[15][36] , \cache_data[15][35] , \cache_data[15][34] ,
         \cache_data[15][33] , \cache_data[15][32] , \cache_data[15][31] ,
         \cache_data[15][30] , \cache_data[15][29] , \cache_data[15][28] ,
         \cache_data[15][27] , \cache_data[15][26] , \cache_data[15][25] ,
         \cache_data[15][24] , \cache_data[15][23] , \cache_data[15][22] ,
         \cache_data[15][21] , \cache_data[15][20] , \cache_data[15][19] ,
         \cache_data[15][18] , \cache_data[15][17] , \cache_data[15][16] ,
         \cache_data[15][15] , \cache_data[15][14] , \cache_data[15][13] ,
         \cache_data[15][12] , \cache_data[15][11] , \cache_data[15][10] ,
         \cache_data[15][9] , \cache_data[15][8] , \cache_data[15][7] ,
         \cache_data[15][6] , \cache_data[15][5] , \cache_data[15][4] ,
         \cache_data[15][3] , \cache_data[15][2] , \cache_data[15][1] ,
         \cache_data[15][0] , \cache_data[14][127] , \cache_data[14][126] ,
         \cache_data[14][125] , \cache_data[14][124] , \cache_data[14][123] ,
         \cache_data[14][122] , \cache_data[14][121] , \cache_data[14][120] ,
         \cache_data[14][119] , \cache_data[14][118] , \cache_data[14][117] ,
         \cache_data[14][116] , \cache_data[14][115] , \cache_data[14][114] ,
         \cache_data[14][113] , \cache_data[14][112] , \cache_data[14][111] ,
         \cache_data[14][110] , \cache_data[14][109] , \cache_data[14][108] ,
         \cache_data[14][107] , \cache_data[14][106] , \cache_data[14][105] ,
         \cache_data[14][104] , \cache_data[14][103] , \cache_data[14][102] ,
         \cache_data[14][101] , \cache_data[14][100] , \cache_data[14][99] ,
         \cache_data[14][98] , \cache_data[14][97] , \cache_data[14][96] ,
         \cache_data[14][95] , \cache_data[14][94] , \cache_data[14][93] ,
         \cache_data[14][92] , \cache_data[14][91] , \cache_data[14][90] ,
         \cache_data[14][89] , \cache_data[14][88] , \cache_data[14][87] ,
         \cache_data[14][86] , \cache_data[14][85] , \cache_data[14][84] ,
         \cache_data[14][83] , \cache_data[14][82] , \cache_data[14][81] ,
         \cache_data[14][80] , \cache_data[14][79] , \cache_data[14][78] ,
         \cache_data[14][77] , \cache_data[14][76] , \cache_data[14][75] ,
         \cache_data[14][74] , \cache_data[14][73] , \cache_data[14][72] ,
         \cache_data[14][71] , \cache_data[14][70] , \cache_data[14][69] ,
         \cache_data[14][68] , \cache_data[14][67] , \cache_data[14][66] ,
         \cache_data[14][65] , \cache_data[14][64] , \cache_data[14][63] ,
         \cache_data[14][62] , \cache_data[14][61] , \cache_data[14][60] ,
         \cache_data[14][59] , \cache_data[14][58] , \cache_data[14][57] ,
         \cache_data[14][56] , \cache_data[14][55] , \cache_data[14][54] ,
         \cache_data[14][53] , \cache_data[14][52] , \cache_data[14][51] ,
         \cache_data[14][50] , \cache_data[14][49] , \cache_data[14][48] ,
         \cache_data[14][47] , \cache_data[14][46] , \cache_data[14][45] ,
         \cache_data[14][44] , \cache_data[14][43] , \cache_data[14][42] ,
         \cache_data[14][41] , \cache_data[14][40] , \cache_data[14][39] ,
         \cache_data[14][38] , \cache_data[14][37] , \cache_data[14][36] ,
         \cache_data[14][35] , \cache_data[14][34] , \cache_data[14][33] ,
         \cache_data[14][32] , \cache_data[14][31] , \cache_data[14][30] ,
         \cache_data[14][29] , \cache_data[14][28] , \cache_data[14][27] ,
         \cache_data[14][26] , \cache_data[14][25] , \cache_data[14][24] ,
         \cache_data[14][23] , \cache_data[14][22] , \cache_data[14][21] ,
         \cache_data[14][20] , \cache_data[14][19] , \cache_data[14][18] ,
         \cache_data[14][17] , \cache_data[14][16] , \cache_data[14][15] ,
         \cache_data[14][14] , \cache_data[14][13] , \cache_data[14][12] ,
         \cache_data[14][11] , \cache_data[14][10] , \cache_data[14][9] ,
         \cache_data[14][8] , \cache_data[14][7] , \cache_data[14][6] ,
         \cache_data[14][5] , \cache_data[14][4] , \cache_data[14][3] ,
         \cache_data[14][2] , \cache_data[14][1] , \cache_data[14][0] ,
         \cache_data[13][127] , \cache_data[13][126] , \cache_data[13][125] ,
         \cache_data[13][124] , \cache_data[13][123] , \cache_data[13][122] ,
         \cache_data[13][121] , \cache_data[13][120] , \cache_data[13][119] ,
         \cache_data[13][118] , \cache_data[13][117] , \cache_data[13][116] ,
         \cache_data[13][115] , \cache_data[13][114] , \cache_data[13][113] ,
         \cache_data[13][112] , \cache_data[13][111] , \cache_data[13][110] ,
         \cache_data[13][109] , \cache_data[13][108] , \cache_data[13][107] ,
         \cache_data[13][106] , \cache_data[13][105] , \cache_data[13][104] ,
         \cache_data[13][103] , \cache_data[13][102] , \cache_data[13][101] ,
         \cache_data[13][100] , \cache_data[13][99] , \cache_data[13][98] ,
         \cache_data[13][97] , \cache_data[13][96] , \cache_data[13][95] ,
         \cache_data[13][94] , \cache_data[13][93] , \cache_data[13][92] ,
         \cache_data[13][91] , \cache_data[13][90] , \cache_data[13][89] ,
         \cache_data[13][88] , \cache_data[13][87] , \cache_data[13][86] ,
         \cache_data[13][85] , \cache_data[13][84] , \cache_data[13][83] ,
         \cache_data[13][82] , \cache_data[13][81] , \cache_data[13][80] ,
         \cache_data[13][79] , \cache_data[13][78] , \cache_data[13][77] ,
         \cache_data[13][76] , \cache_data[13][75] , \cache_data[13][74] ,
         \cache_data[13][73] , \cache_data[13][72] , \cache_data[13][71] ,
         \cache_data[13][70] , \cache_data[13][69] , \cache_data[13][68] ,
         \cache_data[13][67] , \cache_data[13][66] , \cache_data[13][65] ,
         \cache_data[13][64] , \cache_data[13][63] , \cache_data[13][62] ,
         \cache_data[13][61] , \cache_data[13][60] , \cache_data[13][59] ,
         \cache_data[13][58] , \cache_data[13][57] , \cache_data[13][56] ,
         \cache_data[13][55] , \cache_data[13][54] , \cache_data[13][53] ,
         \cache_data[13][52] , \cache_data[13][51] , \cache_data[13][50] ,
         \cache_data[13][49] , \cache_data[13][48] , \cache_data[13][47] ,
         \cache_data[13][46] , \cache_data[13][45] , \cache_data[13][44] ,
         \cache_data[13][43] , \cache_data[13][42] , \cache_data[13][41] ,
         \cache_data[13][40] , \cache_data[13][39] , \cache_data[13][38] ,
         \cache_data[13][37] , \cache_data[13][36] , \cache_data[13][35] ,
         \cache_data[13][34] , \cache_data[13][33] , \cache_data[13][32] ,
         \cache_data[13][31] , \cache_data[13][30] , \cache_data[13][29] ,
         \cache_data[13][28] , \cache_data[13][27] , \cache_data[13][26] ,
         \cache_data[13][25] , \cache_data[13][24] , \cache_data[13][23] ,
         \cache_data[13][22] , \cache_data[13][21] , \cache_data[13][20] ,
         \cache_data[13][19] , \cache_data[13][18] , \cache_data[13][17] ,
         \cache_data[13][16] , \cache_data[13][15] , \cache_data[13][14] ,
         \cache_data[13][13] , \cache_data[13][12] , \cache_data[13][11] ,
         \cache_data[13][10] , \cache_data[13][9] , \cache_data[13][8] ,
         \cache_data[13][7] , \cache_data[13][6] , \cache_data[13][5] ,
         \cache_data[13][4] , \cache_data[13][3] , \cache_data[13][2] ,
         \cache_data[13][1] , \cache_data[13][0] , \cache_data[12][127] ,
         \cache_data[12][126] , \cache_data[12][125] , \cache_data[12][124] ,
         \cache_data[12][123] , \cache_data[12][122] , \cache_data[12][121] ,
         \cache_data[12][120] , \cache_data[12][119] , \cache_data[12][118] ,
         \cache_data[12][117] , \cache_data[12][116] , \cache_data[12][115] ,
         \cache_data[12][114] , \cache_data[12][113] , \cache_data[12][112] ,
         \cache_data[12][111] , \cache_data[12][110] , \cache_data[12][109] ,
         \cache_data[12][108] , \cache_data[12][107] , \cache_data[12][106] ,
         \cache_data[12][105] , \cache_data[12][104] , \cache_data[12][103] ,
         \cache_data[12][102] , \cache_data[12][101] , \cache_data[12][100] ,
         \cache_data[12][99] , \cache_data[12][98] , \cache_data[12][97] ,
         \cache_data[12][96] , \cache_data[12][95] , \cache_data[12][94] ,
         \cache_data[12][93] , \cache_data[12][92] , \cache_data[12][91] ,
         \cache_data[12][90] , \cache_data[12][89] , \cache_data[12][88] ,
         \cache_data[12][87] , \cache_data[12][86] , \cache_data[12][85] ,
         \cache_data[12][84] , \cache_data[12][83] , \cache_data[12][82] ,
         \cache_data[12][81] , \cache_data[12][80] , \cache_data[12][79] ,
         \cache_data[12][78] , \cache_data[12][77] , \cache_data[12][76] ,
         \cache_data[12][75] , \cache_data[12][74] , \cache_data[12][73] ,
         \cache_data[12][72] , \cache_data[12][71] , \cache_data[12][70] ,
         \cache_data[12][69] , \cache_data[12][68] , \cache_data[12][67] ,
         \cache_data[12][66] , \cache_data[12][65] , \cache_data[12][64] ,
         \cache_data[12][63] , \cache_data[12][62] , \cache_data[12][61] ,
         \cache_data[12][60] , \cache_data[12][59] , \cache_data[12][58] ,
         \cache_data[12][57] , \cache_data[12][56] , \cache_data[12][55] ,
         \cache_data[12][54] , \cache_data[12][53] , \cache_data[12][52] ,
         \cache_data[12][51] , \cache_data[12][50] , \cache_data[12][49] ,
         \cache_data[12][48] , \cache_data[12][47] , \cache_data[12][46] ,
         \cache_data[12][45] , \cache_data[12][44] , \cache_data[12][43] ,
         \cache_data[12][42] , \cache_data[12][41] , \cache_data[12][40] ,
         \cache_data[12][39] , \cache_data[12][38] , \cache_data[12][37] ,
         \cache_data[12][36] , \cache_data[12][35] , \cache_data[12][34] ,
         \cache_data[12][33] , \cache_data[12][32] , \cache_data[12][31] ,
         \cache_data[12][30] , \cache_data[12][29] , \cache_data[12][28] ,
         \cache_data[12][27] , \cache_data[12][26] , \cache_data[12][25] ,
         \cache_data[12][24] , \cache_data[12][23] , \cache_data[12][22] ,
         \cache_data[12][21] , \cache_data[12][20] , \cache_data[12][19] ,
         \cache_data[12][18] , \cache_data[12][17] , \cache_data[12][16] ,
         \cache_data[12][15] , \cache_data[12][14] , \cache_data[12][13] ,
         \cache_data[12][12] , \cache_data[12][11] , \cache_data[12][10] ,
         \cache_data[12][9] , \cache_data[12][8] , \cache_data[12][7] ,
         \cache_data[12][6] , \cache_data[12][5] , \cache_data[12][4] ,
         \cache_data[12][3] , \cache_data[12][2] , \cache_data[12][1] ,
         \cache_data[12][0] , \cache_data[11][127] , \cache_data[11][126] ,
         \cache_data[11][125] , \cache_data[11][124] , \cache_data[11][123] ,
         \cache_data[11][122] , \cache_data[11][121] , \cache_data[11][120] ,
         \cache_data[11][119] , \cache_data[11][118] , \cache_data[11][117] ,
         \cache_data[11][116] , \cache_data[11][115] , \cache_data[11][114] ,
         \cache_data[11][113] , \cache_data[11][112] , \cache_data[11][111] ,
         \cache_data[11][110] , \cache_data[11][109] , \cache_data[11][108] ,
         \cache_data[11][107] , \cache_data[11][106] , \cache_data[11][105] ,
         \cache_data[11][104] , \cache_data[11][103] , \cache_data[11][102] ,
         \cache_data[11][101] , \cache_data[11][100] , \cache_data[11][99] ,
         \cache_data[11][98] , \cache_data[11][97] , \cache_data[11][96] ,
         \cache_data[11][95] , \cache_data[11][94] , \cache_data[11][93] ,
         \cache_data[11][92] , \cache_data[11][91] , \cache_data[11][90] ,
         \cache_data[11][89] , \cache_data[11][88] , \cache_data[11][87] ,
         \cache_data[11][86] , \cache_data[11][85] , \cache_data[11][84] ,
         \cache_data[11][83] , \cache_data[11][82] , \cache_data[11][81] ,
         \cache_data[11][80] , \cache_data[11][79] , \cache_data[11][78] ,
         \cache_data[11][77] , \cache_data[11][76] , \cache_data[11][75] ,
         \cache_data[11][74] , \cache_data[11][73] , \cache_data[11][72] ,
         \cache_data[11][71] , \cache_data[11][70] , \cache_data[11][69] ,
         \cache_data[11][68] , \cache_data[11][67] , \cache_data[11][66] ,
         \cache_data[11][65] , \cache_data[11][64] , \cache_data[11][63] ,
         \cache_data[11][62] , \cache_data[11][61] , \cache_data[11][60] ,
         \cache_data[11][59] , \cache_data[11][58] , \cache_data[11][57] ,
         \cache_data[11][56] , \cache_data[11][55] , \cache_data[11][54] ,
         \cache_data[11][53] , \cache_data[11][52] , \cache_data[11][51] ,
         \cache_data[11][50] , \cache_data[11][49] , \cache_data[11][48] ,
         \cache_data[11][47] , \cache_data[11][46] , \cache_data[11][45] ,
         \cache_data[11][44] , \cache_data[11][43] , \cache_data[11][42] ,
         \cache_data[11][41] , \cache_data[11][40] , \cache_data[11][39] ,
         \cache_data[11][38] , \cache_data[11][37] , \cache_data[11][36] ,
         \cache_data[11][35] , \cache_data[11][34] , \cache_data[11][33] ,
         \cache_data[11][32] , \cache_data[11][31] , \cache_data[11][30] ,
         \cache_data[11][29] , \cache_data[11][28] , \cache_data[11][27] ,
         \cache_data[11][26] , \cache_data[11][25] , \cache_data[11][24] ,
         \cache_data[11][23] , \cache_data[11][22] , \cache_data[11][21] ,
         \cache_data[11][20] , \cache_data[11][19] , \cache_data[11][18] ,
         \cache_data[11][17] , \cache_data[11][16] , \cache_data[11][15] ,
         \cache_data[11][14] , \cache_data[11][13] , \cache_data[11][12] ,
         \cache_data[11][11] , \cache_data[11][10] , \cache_data[11][9] ,
         \cache_data[11][8] , \cache_data[11][7] , \cache_data[11][6] ,
         \cache_data[11][5] , \cache_data[11][4] , \cache_data[11][3] ,
         \cache_data[11][2] , \cache_data[11][1] , \cache_data[11][0] ,
         \cache_data[10][127] , \cache_data[10][126] , \cache_data[10][125] ,
         \cache_data[10][124] , \cache_data[10][123] , \cache_data[10][122] ,
         \cache_data[10][121] , \cache_data[10][120] , \cache_data[10][119] ,
         \cache_data[10][118] , \cache_data[10][117] , \cache_data[10][116] ,
         \cache_data[10][115] , \cache_data[10][114] , \cache_data[10][113] ,
         \cache_data[10][112] , \cache_data[10][111] , \cache_data[10][110] ,
         \cache_data[10][109] , \cache_data[10][108] , \cache_data[10][107] ,
         \cache_data[10][106] , \cache_data[10][105] , \cache_data[10][104] ,
         \cache_data[10][103] , \cache_data[10][102] , \cache_data[10][101] ,
         \cache_data[10][100] , \cache_data[10][99] , \cache_data[10][98] ,
         \cache_data[10][97] , \cache_data[10][96] , \cache_data[10][95] ,
         \cache_data[10][94] , \cache_data[10][93] , \cache_data[10][92] ,
         \cache_data[10][91] , \cache_data[10][90] , \cache_data[10][89] ,
         \cache_data[10][88] , \cache_data[10][87] , \cache_data[10][86] ,
         \cache_data[10][85] , \cache_data[10][84] , \cache_data[10][83] ,
         \cache_data[10][82] , \cache_data[10][81] , \cache_data[10][80] ,
         \cache_data[10][79] , \cache_data[10][78] , \cache_data[10][77] ,
         \cache_data[10][76] , \cache_data[10][75] , \cache_data[10][74] ,
         \cache_data[10][73] , \cache_data[10][72] , \cache_data[10][71] ,
         \cache_data[10][70] , \cache_data[10][69] , \cache_data[10][68] ,
         \cache_data[10][67] , \cache_data[10][66] , \cache_data[10][65] ,
         \cache_data[10][64] , \cache_data[10][63] , \cache_data[10][62] ,
         \cache_data[10][61] , \cache_data[10][60] , \cache_data[10][59] ,
         \cache_data[10][58] , \cache_data[10][57] , \cache_data[10][56] ,
         \cache_data[10][55] , \cache_data[10][54] , \cache_data[10][53] ,
         \cache_data[10][52] , \cache_data[10][51] , \cache_data[10][50] ,
         \cache_data[10][49] , \cache_data[10][48] , \cache_data[10][47] ,
         \cache_data[10][46] , \cache_data[10][45] , \cache_data[10][44] ,
         \cache_data[10][43] , \cache_data[10][42] , \cache_data[10][41] ,
         \cache_data[10][40] , \cache_data[10][39] , \cache_data[10][38] ,
         \cache_data[10][37] , \cache_data[10][36] , \cache_data[10][35] ,
         \cache_data[10][34] , \cache_data[10][33] , \cache_data[10][32] ,
         \cache_data[10][31] , \cache_data[10][30] , \cache_data[10][29] ,
         \cache_data[10][28] , \cache_data[10][27] , \cache_data[10][26] ,
         \cache_data[10][25] , \cache_data[10][24] , \cache_data[10][23] ,
         \cache_data[10][22] , \cache_data[10][21] , \cache_data[10][20] ,
         \cache_data[10][19] , \cache_data[10][18] , \cache_data[10][17] ,
         \cache_data[10][16] , \cache_data[10][15] , \cache_data[10][14] ,
         \cache_data[10][13] , \cache_data[10][12] , \cache_data[10][11] ,
         \cache_data[10][10] , \cache_data[10][9] , \cache_data[10][8] ,
         \cache_data[10][7] , \cache_data[10][6] , \cache_data[10][5] ,
         \cache_data[10][4] , \cache_data[10][3] , \cache_data[10][2] ,
         \cache_data[10][1] , \cache_data[10][0] , \cache_data[9][127] ,
         \cache_data[9][126] , \cache_data[9][125] , \cache_data[9][124] ,
         \cache_data[9][123] , \cache_data[9][122] , \cache_data[9][121] ,
         \cache_data[9][120] , \cache_data[9][119] , \cache_data[9][118] ,
         \cache_data[9][117] , \cache_data[9][116] , \cache_data[9][115] ,
         \cache_data[9][114] , \cache_data[9][113] , \cache_data[9][112] ,
         \cache_data[9][111] , \cache_data[9][110] , \cache_data[9][109] ,
         \cache_data[9][108] , \cache_data[9][107] , \cache_data[9][106] ,
         \cache_data[9][105] , \cache_data[9][104] , \cache_data[9][103] ,
         \cache_data[9][102] , \cache_data[9][101] , \cache_data[9][100] ,
         \cache_data[9][99] , \cache_data[9][98] , \cache_data[9][97] ,
         \cache_data[9][96] , \cache_data[9][95] , \cache_data[9][94] ,
         \cache_data[9][93] , \cache_data[9][92] , \cache_data[9][91] ,
         \cache_data[9][90] , \cache_data[9][89] , \cache_data[9][88] ,
         \cache_data[9][87] , \cache_data[9][86] , \cache_data[9][85] ,
         \cache_data[9][84] , \cache_data[9][83] , \cache_data[9][82] ,
         \cache_data[9][81] , \cache_data[9][80] , \cache_data[9][79] ,
         \cache_data[9][78] , \cache_data[9][77] , \cache_data[9][76] ,
         \cache_data[9][75] , \cache_data[9][74] , \cache_data[9][73] ,
         \cache_data[9][72] , \cache_data[9][71] , \cache_data[9][70] ,
         \cache_data[9][69] , \cache_data[9][68] , \cache_data[9][67] ,
         \cache_data[9][66] , \cache_data[9][65] , \cache_data[9][64] ,
         \cache_data[9][63] , \cache_data[9][62] , \cache_data[9][61] ,
         \cache_data[9][60] , \cache_data[9][59] , \cache_data[9][58] ,
         \cache_data[9][57] , \cache_data[9][56] , \cache_data[9][55] ,
         \cache_data[9][54] , \cache_data[9][53] , \cache_data[9][52] ,
         \cache_data[9][51] , \cache_data[9][50] , \cache_data[9][49] ,
         \cache_data[9][48] , \cache_data[9][47] , \cache_data[9][46] ,
         \cache_data[9][45] , \cache_data[9][44] , \cache_data[9][43] ,
         \cache_data[9][42] , \cache_data[9][41] , \cache_data[9][40] ,
         \cache_data[9][39] , \cache_data[9][38] , \cache_data[9][37] ,
         \cache_data[9][36] , \cache_data[9][35] , \cache_data[9][34] ,
         \cache_data[9][33] , \cache_data[9][32] , \cache_data[9][31] ,
         \cache_data[9][30] , \cache_data[9][29] , \cache_data[9][28] ,
         \cache_data[9][27] , \cache_data[9][26] , \cache_data[9][25] ,
         \cache_data[9][24] , \cache_data[9][23] , \cache_data[9][22] ,
         \cache_data[9][21] , \cache_data[9][20] , \cache_data[9][19] ,
         \cache_data[9][18] , \cache_data[9][17] , \cache_data[9][16] ,
         \cache_data[9][15] , \cache_data[9][14] , \cache_data[9][13] ,
         \cache_data[9][12] , \cache_data[9][11] , \cache_data[9][10] ,
         \cache_data[9][9] , \cache_data[9][8] , \cache_data[9][7] ,
         \cache_data[9][6] , \cache_data[9][5] , \cache_data[9][4] ,
         \cache_data[9][3] , \cache_data[9][2] , \cache_data[9][1] ,
         \cache_data[9][0] , \cache_data[8][127] , \cache_data[8][126] ,
         \cache_data[8][125] , \cache_data[8][124] , \cache_data[8][123] ,
         \cache_data[8][122] , \cache_data[8][121] , \cache_data[8][120] ,
         \cache_data[8][119] , \cache_data[8][118] , \cache_data[8][117] ,
         \cache_data[8][116] , \cache_data[8][115] , \cache_data[8][114] ,
         \cache_data[8][113] , \cache_data[8][112] , \cache_data[8][111] ,
         \cache_data[8][110] , \cache_data[8][109] , \cache_data[8][108] ,
         \cache_data[8][107] , \cache_data[8][106] , \cache_data[8][105] ,
         \cache_data[8][104] , \cache_data[8][103] , \cache_data[8][102] ,
         \cache_data[8][101] , \cache_data[8][100] , \cache_data[8][99] ,
         \cache_data[8][98] , \cache_data[8][97] , \cache_data[8][96] ,
         \cache_data[8][95] , \cache_data[8][94] , \cache_data[8][93] ,
         \cache_data[8][92] , \cache_data[8][91] , \cache_data[8][90] ,
         \cache_data[8][89] , \cache_data[8][88] , \cache_data[8][87] ,
         \cache_data[8][86] , \cache_data[8][85] , \cache_data[8][84] ,
         \cache_data[8][83] , \cache_data[8][82] , \cache_data[8][81] ,
         \cache_data[8][80] , \cache_data[8][79] , \cache_data[8][78] ,
         \cache_data[8][77] , \cache_data[8][76] , \cache_data[8][75] ,
         \cache_data[8][74] , \cache_data[8][73] , \cache_data[8][72] ,
         \cache_data[8][71] , \cache_data[8][70] , \cache_data[8][69] ,
         \cache_data[8][68] , \cache_data[8][67] , \cache_data[8][66] ,
         \cache_data[8][65] , \cache_data[8][64] , \cache_data[8][63] ,
         \cache_data[8][62] , \cache_data[8][61] , \cache_data[8][60] ,
         \cache_data[8][59] , \cache_data[8][58] , \cache_data[8][57] ,
         \cache_data[8][56] , \cache_data[8][55] , \cache_data[8][54] ,
         \cache_data[8][53] , \cache_data[8][52] , \cache_data[8][51] ,
         \cache_data[8][50] , \cache_data[8][49] , \cache_data[8][48] ,
         \cache_data[8][47] , \cache_data[8][46] , \cache_data[8][45] ,
         \cache_data[8][44] , \cache_data[8][43] , \cache_data[8][42] ,
         \cache_data[8][41] , \cache_data[8][40] , \cache_data[8][39] ,
         \cache_data[8][38] , \cache_data[8][37] , \cache_data[8][36] ,
         \cache_data[8][35] , \cache_data[8][34] , \cache_data[8][33] ,
         \cache_data[8][32] , \cache_data[8][31] , \cache_data[8][30] ,
         \cache_data[8][29] , \cache_data[8][28] , \cache_data[8][27] ,
         \cache_data[8][26] , \cache_data[8][25] , \cache_data[8][24] ,
         \cache_data[8][23] , \cache_data[8][22] , \cache_data[8][21] ,
         \cache_data[8][20] , \cache_data[8][19] , \cache_data[8][18] ,
         \cache_data[8][17] , \cache_data[8][16] , \cache_data[8][15] ,
         \cache_data[8][14] , \cache_data[8][13] , \cache_data[8][12] ,
         \cache_data[8][11] , \cache_data[8][10] , \cache_data[8][9] ,
         \cache_data[8][8] , \cache_data[8][7] , \cache_data[8][6] ,
         \cache_data[8][5] , \cache_data[8][4] , \cache_data[8][3] ,
         \cache_data[8][2] , \cache_data[8][1] , \cache_data[8][0] ,
         \cache_data[7][127] , \cache_data[7][126] , \cache_data[7][125] ,
         \cache_data[7][124] , \cache_data[7][123] , \cache_data[7][122] ,
         \cache_data[7][121] , \cache_data[7][120] , \cache_data[7][119] ,
         \cache_data[7][118] , \cache_data[7][117] , \cache_data[7][116] ,
         \cache_data[7][115] , \cache_data[7][114] , \cache_data[7][113] ,
         \cache_data[7][112] , \cache_data[7][111] , \cache_data[7][110] ,
         \cache_data[7][109] , \cache_data[7][108] , \cache_data[7][107] ,
         \cache_data[7][106] , \cache_data[7][105] , \cache_data[7][104] ,
         \cache_data[7][103] , \cache_data[7][102] , \cache_data[7][101] ,
         \cache_data[7][100] , \cache_data[7][99] , \cache_data[7][98] ,
         \cache_data[7][97] , \cache_data[7][96] , \cache_data[7][95] ,
         \cache_data[7][94] , \cache_data[7][93] , \cache_data[7][92] ,
         \cache_data[7][91] , \cache_data[7][90] , \cache_data[7][89] ,
         \cache_data[7][88] , \cache_data[7][87] , \cache_data[7][86] ,
         \cache_data[7][85] , \cache_data[7][84] , \cache_data[7][83] ,
         \cache_data[7][82] , \cache_data[7][81] , \cache_data[7][80] ,
         \cache_data[7][79] , \cache_data[7][78] , \cache_data[7][77] ,
         \cache_data[7][76] , \cache_data[7][75] , \cache_data[7][74] ,
         \cache_data[7][73] , \cache_data[7][72] , \cache_data[7][71] ,
         \cache_data[7][70] , \cache_data[7][69] , \cache_data[7][68] ,
         \cache_data[7][67] , \cache_data[7][66] , \cache_data[7][65] ,
         \cache_data[7][64] , \cache_data[7][63] , \cache_data[7][62] ,
         \cache_data[7][61] , \cache_data[7][60] , \cache_data[7][59] ,
         \cache_data[7][58] , \cache_data[7][57] , \cache_data[7][56] ,
         \cache_data[7][55] , \cache_data[7][54] , \cache_data[7][53] ,
         \cache_data[7][52] , \cache_data[7][51] , \cache_data[7][50] ,
         \cache_data[7][49] , \cache_data[7][48] , \cache_data[7][47] ,
         \cache_data[7][46] , \cache_data[7][45] , \cache_data[7][44] ,
         \cache_data[7][43] , \cache_data[7][42] , \cache_data[7][41] ,
         \cache_data[7][40] , \cache_data[7][39] , \cache_data[7][38] ,
         \cache_data[7][37] , \cache_data[7][36] , \cache_data[7][35] ,
         \cache_data[7][34] , \cache_data[7][33] , \cache_data[7][32] ,
         \cache_data[7][31] , \cache_data[7][30] , \cache_data[7][29] ,
         \cache_data[7][28] , \cache_data[7][27] , \cache_data[7][26] ,
         \cache_data[7][25] , \cache_data[7][24] , \cache_data[7][23] ,
         \cache_data[7][22] , \cache_data[7][21] , \cache_data[7][20] ,
         \cache_data[7][19] , \cache_data[7][18] , \cache_data[7][17] ,
         \cache_data[7][16] , \cache_data[7][15] , \cache_data[7][14] ,
         \cache_data[7][13] , \cache_data[7][12] , \cache_data[7][11] ,
         \cache_data[7][10] , \cache_data[7][9] , \cache_data[7][8] ,
         \cache_data[7][7] , \cache_data[7][6] , \cache_data[7][5] ,
         \cache_data[7][4] , \cache_data[7][3] , \cache_data[7][2] ,
         \cache_data[7][1] , \cache_data[7][0] , \cache_data[6][127] ,
         \cache_data[6][126] , \cache_data[6][125] , \cache_data[6][124] ,
         \cache_data[6][123] , \cache_data[6][122] , \cache_data[6][121] ,
         \cache_data[6][120] , \cache_data[6][119] , \cache_data[6][118] ,
         \cache_data[6][117] , \cache_data[6][116] , \cache_data[6][115] ,
         \cache_data[6][114] , \cache_data[6][113] , \cache_data[6][112] ,
         \cache_data[6][111] , \cache_data[6][110] , \cache_data[6][109] ,
         \cache_data[6][108] , \cache_data[6][107] , \cache_data[6][106] ,
         \cache_data[6][105] , \cache_data[6][104] , \cache_data[6][103] ,
         \cache_data[6][102] , \cache_data[6][101] , \cache_data[6][100] ,
         \cache_data[6][99] , \cache_data[6][98] , \cache_data[6][97] ,
         \cache_data[6][96] , \cache_data[6][95] , \cache_data[6][94] ,
         \cache_data[6][93] , \cache_data[6][92] , \cache_data[6][91] ,
         \cache_data[6][90] , \cache_data[6][89] , \cache_data[6][88] ,
         \cache_data[6][87] , \cache_data[6][86] , \cache_data[6][85] ,
         \cache_data[6][84] , \cache_data[6][83] , \cache_data[6][82] ,
         \cache_data[6][81] , \cache_data[6][80] , \cache_data[6][79] ,
         \cache_data[6][78] , \cache_data[6][77] , \cache_data[6][76] ,
         \cache_data[6][75] , \cache_data[6][74] , \cache_data[6][73] ,
         \cache_data[6][72] , \cache_data[6][71] , \cache_data[6][70] ,
         \cache_data[6][69] , \cache_data[6][68] , \cache_data[6][67] ,
         \cache_data[6][66] , \cache_data[6][65] , \cache_data[6][64] ,
         \cache_data[6][63] , \cache_data[6][62] , \cache_data[6][61] ,
         \cache_data[6][60] , \cache_data[6][59] , \cache_data[6][58] ,
         \cache_data[6][57] , \cache_data[6][56] , \cache_data[6][55] ,
         \cache_data[6][54] , \cache_data[6][53] , \cache_data[6][52] ,
         \cache_data[6][51] , \cache_data[6][50] , \cache_data[6][49] ,
         \cache_data[6][48] , \cache_data[6][47] , \cache_data[6][46] ,
         \cache_data[6][45] , \cache_data[6][44] , \cache_data[6][43] ,
         \cache_data[6][42] , \cache_data[6][41] , \cache_data[6][40] ,
         \cache_data[6][39] , \cache_data[6][38] , \cache_data[6][37] ,
         \cache_data[6][36] , \cache_data[6][35] , \cache_data[6][34] ,
         \cache_data[6][33] , \cache_data[6][32] , \cache_data[6][31] ,
         \cache_data[6][30] , \cache_data[6][29] , \cache_data[6][28] ,
         \cache_data[6][27] , \cache_data[6][26] , \cache_data[6][25] ,
         \cache_data[6][24] , \cache_data[6][23] , \cache_data[6][22] ,
         \cache_data[6][21] , \cache_data[6][20] , \cache_data[6][19] ,
         \cache_data[6][18] , \cache_data[6][17] , \cache_data[6][16] ,
         \cache_data[6][15] , \cache_data[6][14] , \cache_data[6][13] ,
         \cache_data[6][12] , \cache_data[6][11] , \cache_data[6][10] ,
         \cache_data[6][9] , \cache_data[6][8] , \cache_data[6][7] ,
         \cache_data[6][6] , \cache_data[6][5] , \cache_data[6][4] ,
         \cache_data[6][3] , \cache_data[6][2] , \cache_data[6][1] ,
         \cache_data[6][0] , \cache_data[5][127] , \cache_data[5][126] ,
         \cache_data[5][125] , \cache_data[5][124] , \cache_data[5][123] ,
         \cache_data[5][122] , \cache_data[5][121] , \cache_data[5][120] ,
         \cache_data[5][119] , \cache_data[5][118] , \cache_data[5][117] ,
         \cache_data[5][116] , \cache_data[5][115] , \cache_data[5][114] ,
         \cache_data[5][113] , \cache_data[5][112] , \cache_data[5][111] ,
         \cache_data[5][110] , \cache_data[5][109] , \cache_data[5][108] ,
         \cache_data[5][107] , \cache_data[5][106] , \cache_data[5][105] ,
         \cache_data[5][104] , \cache_data[5][103] , \cache_data[5][102] ,
         \cache_data[5][101] , \cache_data[5][100] , \cache_data[5][99] ,
         \cache_data[5][98] , \cache_data[5][97] , \cache_data[5][96] ,
         \cache_data[5][95] , \cache_data[5][94] , \cache_data[5][93] ,
         \cache_data[5][92] , \cache_data[5][91] , \cache_data[5][90] ,
         \cache_data[5][89] , \cache_data[5][88] , \cache_data[5][87] ,
         \cache_data[5][86] , \cache_data[5][85] , \cache_data[5][84] ,
         \cache_data[5][83] , \cache_data[5][82] , \cache_data[5][81] ,
         \cache_data[5][80] , \cache_data[5][79] , \cache_data[5][78] ,
         \cache_data[5][77] , \cache_data[5][76] , \cache_data[5][75] ,
         \cache_data[5][74] , \cache_data[5][73] , \cache_data[5][72] ,
         \cache_data[5][71] , \cache_data[5][70] , \cache_data[5][69] ,
         \cache_data[5][68] , \cache_data[5][67] , \cache_data[5][66] ,
         \cache_data[5][65] , \cache_data[5][64] , \cache_data[5][63] ,
         \cache_data[5][62] , \cache_data[5][61] , \cache_data[5][60] ,
         \cache_data[5][59] , \cache_data[5][58] , \cache_data[5][57] ,
         \cache_data[5][56] , \cache_data[5][55] , \cache_data[5][54] ,
         \cache_data[5][53] , \cache_data[5][52] , \cache_data[5][51] ,
         \cache_data[5][50] , \cache_data[5][49] , \cache_data[5][48] ,
         \cache_data[5][47] , \cache_data[5][46] , \cache_data[5][45] ,
         \cache_data[5][44] , \cache_data[5][43] , \cache_data[5][42] ,
         \cache_data[5][41] , \cache_data[5][40] , \cache_data[5][39] ,
         \cache_data[5][38] , \cache_data[5][37] , \cache_data[5][36] ,
         \cache_data[5][35] , \cache_data[5][34] , \cache_data[5][33] ,
         \cache_data[5][32] , \cache_data[5][31] , \cache_data[5][30] ,
         \cache_data[5][29] , \cache_data[5][28] , \cache_data[5][27] ,
         \cache_data[5][26] , \cache_data[5][25] , \cache_data[5][24] ,
         \cache_data[5][23] , \cache_data[5][22] , \cache_data[5][21] ,
         \cache_data[5][20] , \cache_data[5][19] , \cache_data[5][18] ,
         \cache_data[5][17] , \cache_data[5][16] , \cache_data[5][15] ,
         \cache_data[5][14] , \cache_data[5][13] , \cache_data[5][12] ,
         \cache_data[5][11] , \cache_data[5][10] , \cache_data[5][9] ,
         \cache_data[5][8] , \cache_data[5][7] , \cache_data[5][6] ,
         \cache_data[5][5] , \cache_data[5][4] , \cache_data[5][3] ,
         \cache_data[5][2] , \cache_data[5][1] , \cache_data[5][0] ,
         \cache_data[4][127] , \cache_data[4][126] , \cache_data[4][125] ,
         \cache_data[4][124] , \cache_data[4][123] , \cache_data[4][122] ,
         \cache_data[4][121] , \cache_data[4][120] , \cache_data[4][119] ,
         \cache_data[4][118] , \cache_data[4][117] , \cache_data[4][116] ,
         \cache_data[4][115] , \cache_data[4][114] , \cache_data[4][113] ,
         \cache_data[4][112] , \cache_data[4][111] , \cache_data[4][110] ,
         \cache_data[4][109] , \cache_data[4][108] , \cache_data[4][107] ,
         \cache_data[4][106] , \cache_data[4][105] , \cache_data[4][104] ,
         \cache_data[4][103] , \cache_data[4][102] , \cache_data[4][101] ,
         \cache_data[4][100] , \cache_data[4][99] , \cache_data[4][98] ,
         \cache_data[4][97] , \cache_data[4][96] , \cache_data[4][95] ,
         \cache_data[4][94] , \cache_data[4][93] , \cache_data[4][92] ,
         \cache_data[4][91] , \cache_data[4][90] , \cache_data[4][89] ,
         \cache_data[4][88] , \cache_data[4][87] , \cache_data[4][86] ,
         \cache_data[4][85] , \cache_data[4][84] , \cache_data[4][83] ,
         \cache_data[4][82] , \cache_data[4][81] , \cache_data[4][80] ,
         \cache_data[4][79] , \cache_data[4][78] , \cache_data[4][77] ,
         \cache_data[4][76] , \cache_data[4][75] , \cache_data[4][74] ,
         \cache_data[4][73] , \cache_data[4][72] , \cache_data[4][71] ,
         \cache_data[4][70] , \cache_data[4][69] , \cache_data[4][68] ,
         \cache_data[4][67] , \cache_data[4][66] , \cache_data[4][65] ,
         \cache_data[4][64] , \cache_data[4][63] , \cache_data[4][62] ,
         \cache_data[4][61] , \cache_data[4][60] , \cache_data[4][59] ,
         \cache_data[4][58] , \cache_data[4][57] , \cache_data[4][56] ,
         \cache_data[4][55] , \cache_data[4][54] , \cache_data[4][53] ,
         \cache_data[4][52] , \cache_data[4][51] , \cache_data[4][50] ,
         \cache_data[4][49] , \cache_data[4][48] , \cache_data[4][47] ,
         \cache_data[4][46] , \cache_data[4][45] , \cache_data[4][44] ,
         \cache_data[4][43] , \cache_data[4][42] , \cache_data[4][41] ,
         \cache_data[4][40] , \cache_data[4][39] , \cache_data[4][38] ,
         \cache_data[4][37] , \cache_data[4][36] , \cache_data[4][35] ,
         \cache_data[4][34] , \cache_data[4][33] , \cache_data[4][32] ,
         \cache_data[4][31] , \cache_data[4][30] , \cache_data[4][29] ,
         \cache_data[4][28] , \cache_data[4][27] , \cache_data[4][26] ,
         \cache_data[4][25] , \cache_data[4][24] , \cache_data[4][23] ,
         \cache_data[4][22] , \cache_data[4][21] , \cache_data[4][20] ,
         \cache_data[4][19] , \cache_data[4][18] , \cache_data[4][17] ,
         \cache_data[4][16] , \cache_data[4][15] , \cache_data[4][14] ,
         \cache_data[4][13] , \cache_data[4][12] , \cache_data[4][11] ,
         \cache_data[4][10] , \cache_data[4][9] , \cache_data[4][8] ,
         \cache_data[4][7] , \cache_data[4][6] , \cache_data[4][5] ,
         \cache_data[4][4] , \cache_data[4][3] , \cache_data[4][2] ,
         \cache_data[4][1] , \cache_data[4][0] , \cache_data[3][127] ,
         \cache_data[3][126] , \cache_data[3][125] , \cache_data[3][124] ,
         \cache_data[3][123] , \cache_data[3][122] , \cache_data[3][121] ,
         \cache_data[3][120] , \cache_data[3][119] , \cache_data[3][118] ,
         \cache_data[3][117] , \cache_data[3][116] , \cache_data[3][115] ,
         \cache_data[3][114] , \cache_data[3][113] , \cache_data[3][112] ,
         \cache_data[3][111] , \cache_data[3][110] , \cache_data[3][109] ,
         \cache_data[3][108] , \cache_data[3][107] , \cache_data[3][106] ,
         \cache_data[3][105] , \cache_data[3][104] , \cache_data[3][103] ,
         \cache_data[3][102] , \cache_data[3][101] , \cache_data[3][100] ,
         \cache_data[3][99] , \cache_data[3][98] , \cache_data[3][97] ,
         \cache_data[3][96] , \cache_data[3][95] , \cache_data[3][94] ,
         \cache_data[3][93] , \cache_data[3][92] , \cache_data[3][91] ,
         \cache_data[3][90] , \cache_data[3][89] , \cache_data[3][88] ,
         \cache_data[3][87] , \cache_data[3][86] , \cache_data[3][85] ,
         \cache_data[3][84] , \cache_data[3][83] , \cache_data[3][82] ,
         \cache_data[3][81] , \cache_data[3][80] , \cache_data[3][79] ,
         \cache_data[3][78] , \cache_data[3][77] , \cache_data[3][76] ,
         \cache_data[3][75] , \cache_data[3][74] , \cache_data[3][73] ,
         \cache_data[3][72] , \cache_data[3][71] , \cache_data[3][70] ,
         \cache_data[3][69] , \cache_data[3][68] , \cache_data[3][67] ,
         \cache_data[3][66] , \cache_data[3][65] , \cache_data[3][64] ,
         \cache_data[3][63] , \cache_data[3][62] , \cache_data[3][61] ,
         \cache_data[3][60] , \cache_data[3][59] , \cache_data[3][58] ,
         \cache_data[3][57] , \cache_data[3][56] , \cache_data[3][55] ,
         \cache_data[3][54] , \cache_data[3][53] , \cache_data[3][52] ,
         \cache_data[3][51] , \cache_data[3][50] , \cache_data[3][49] ,
         \cache_data[3][48] , \cache_data[3][47] , \cache_data[3][46] ,
         \cache_data[3][45] , \cache_data[3][44] , \cache_data[3][43] ,
         \cache_data[3][42] , \cache_data[3][41] , \cache_data[3][40] ,
         \cache_data[3][39] , \cache_data[3][38] , \cache_data[3][37] ,
         \cache_data[3][36] , \cache_data[3][35] , \cache_data[3][34] ,
         \cache_data[3][33] , \cache_data[3][32] , \cache_data[3][31] ,
         \cache_data[3][30] , \cache_data[3][29] , \cache_data[3][28] ,
         \cache_data[3][27] , \cache_data[3][26] , \cache_data[3][25] ,
         \cache_data[3][24] , \cache_data[3][23] , \cache_data[3][22] ,
         \cache_data[3][21] , \cache_data[3][20] , \cache_data[3][19] ,
         \cache_data[3][18] , \cache_data[3][17] , \cache_data[3][16] ,
         \cache_data[3][15] , \cache_data[3][14] , \cache_data[3][13] ,
         \cache_data[3][12] , \cache_data[3][11] , \cache_data[3][10] ,
         \cache_data[3][9] , \cache_data[3][8] , \cache_data[3][7] ,
         \cache_data[3][6] , \cache_data[3][5] , \cache_data[3][4] ,
         \cache_data[3][3] , \cache_data[3][2] , \cache_data[3][1] ,
         \cache_data[3][0] , \cache_data[2][127] , \cache_data[2][126] ,
         \cache_data[2][125] , \cache_data[2][124] , \cache_data[2][123] ,
         \cache_data[2][122] , \cache_data[2][121] , \cache_data[2][120] ,
         \cache_data[2][119] , \cache_data[2][118] , \cache_data[2][117] ,
         \cache_data[2][116] , \cache_data[2][115] , \cache_data[2][114] ,
         \cache_data[2][113] , \cache_data[2][112] , \cache_data[2][111] ,
         \cache_data[2][110] , \cache_data[2][109] , \cache_data[2][108] ,
         \cache_data[2][107] , \cache_data[2][106] , \cache_data[2][105] ,
         \cache_data[2][104] , \cache_data[2][103] , \cache_data[2][102] ,
         \cache_data[2][101] , \cache_data[2][100] , \cache_data[2][99] ,
         \cache_data[2][98] , \cache_data[2][97] , \cache_data[2][96] ,
         \cache_data[2][95] , \cache_data[2][94] , \cache_data[2][93] ,
         \cache_data[2][92] , \cache_data[2][91] , \cache_data[2][90] ,
         \cache_data[2][89] , \cache_data[2][88] , \cache_data[2][87] ,
         \cache_data[2][86] , \cache_data[2][85] , \cache_data[2][84] ,
         \cache_data[2][83] , \cache_data[2][82] , \cache_data[2][81] ,
         \cache_data[2][80] , \cache_data[2][79] , \cache_data[2][78] ,
         \cache_data[2][77] , \cache_data[2][76] , \cache_data[2][75] ,
         \cache_data[2][74] , \cache_data[2][73] , \cache_data[2][72] ,
         \cache_data[2][71] , \cache_data[2][70] , \cache_data[2][69] ,
         \cache_data[2][68] , \cache_data[2][67] , \cache_data[2][66] ,
         \cache_data[2][65] , \cache_data[2][64] , \cache_data[2][63] ,
         \cache_data[2][62] , \cache_data[2][61] , \cache_data[2][60] ,
         \cache_data[2][59] , \cache_data[2][58] , \cache_data[2][57] ,
         \cache_data[2][56] , \cache_data[2][55] , \cache_data[2][54] ,
         \cache_data[2][53] , \cache_data[2][52] , \cache_data[2][51] ,
         \cache_data[2][50] , \cache_data[2][49] , \cache_data[2][48] ,
         \cache_data[2][47] , \cache_data[2][46] , \cache_data[2][45] ,
         \cache_data[2][44] , \cache_data[2][43] , \cache_data[2][42] ,
         \cache_data[2][41] , \cache_data[2][40] , \cache_data[2][39] ,
         \cache_data[2][38] , \cache_data[2][37] , \cache_data[2][36] ,
         \cache_data[2][35] , \cache_data[2][34] , \cache_data[2][33] ,
         \cache_data[2][32] , \cache_data[2][31] , \cache_data[2][30] ,
         \cache_data[2][29] , \cache_data[2][28] , \cache_data[2][27] ,
         \cache_data[2][26] , \cache_data[2][25] , \cache_data[2][24] ,
         \cache_data[2][23] , \cache_data[2][22] , \cache_data[2][21] ,
         \cache_data[2][20] , \cache_data[2][19] , \cache_data[2][18] ,
         \cache_data[2][17] , \cache_data[2][16] , \cache_data[2][15] ,
         \cache_data[2][14] , \cache_data[2][13] , \cache_data[2][12] ,
         \cache_data[2][11] , \cache_data[2][10] , \cache_data[2][9] ,
         \cache_data[2][8] , \cache_data[2][7] , \cache_data[2][6] ,
         \cache_data[2][5] , \cache_data[2][4] , \cache_data[2][3] ,
         \cache_data[2][2] , \cache_data[2][1] , \cache_data[2][0] ,
         \cache_data[1][127] , \cache_data[1][126] , \cache_data[1][125] ,
         \cache_data[1][124] , \cache_data[1][123] , \cache_data[1][122] ,
         \cache_data[1][121] , \cache_data[1][120] , \cache_data[1][119] ,
         \cache_data[1][118] , \cache_data[1][117] , \cache_data[1][116] ,
         \cache_data[1][115] , \cache_data[1][114] , \cache_data[1][113] ,
         \cache_data[1][112] , \cache_data[1][111] , \cache_data[1][110] ,
         \cache_data[1][109] , \cache_data[1][108] , \cache_data[1][107] ,
         \cache_data[1][106] , \cache_data[1][105] , \cache_data[1][104] ,
         \cache_data[1][103] , \cache_data[1][102] , \cache_data[1][101] ,
         \cache_data[1][100] , \cache_data[1][99] , \cache_data[1][98] ,
         \cache_data[1][97] , \cache_data[1][96] , \cache_data[1][95] ,
         \cache_data[1][94] , \cache_data[1][93] , \cache_data[1][92] ,
         \cache_data[1][91] , \cache_data[1][90] , \cache_data[1][89] ,
         \cache_data[1][88] , \cache_data[1][87] , \cache_data[1][86] ,
         \cache_data[1][85] , \cache_data[1][84] , \cache_data[1][83] ,
         \cache_data[1][82] , \cache_data[1][81] , \cache_data[1][80] ,
         \cache_data[1][79] , \cache_data[1][78] , \cache_data[1][77] ,
         \cache_data[1][76] , \cache_data[1][75] , \cache_data[1][74] ,
         \cache_data[1][73] , \cache_data[1][72] , \cache_data[1][71] ,
         \cache_data[1][70] , \cache_data[1][69] , \cache_data[1][68] ,
         \cache_data[1][67] , \cache_data[1][66] , \cache_data[1][65] ,
         \cache_data[1][64] , \cache_data[1][63] , \cache_data[1][62] ,
         \cache_data[1][61] , \cache_data[1][60] , \cache_data[1][59] ,
         \cache_data[1][58] , \cache_data[1][57] , \cache_data[1][56] ,
         \cache_data[1][55] , \cache_data[1][54] , \cache_data[1][53] ,
         \cache_data[1][52] , \cache_data[1][51] , \cache_data[1][50] ,
         \cache_data[1][49] , \cache_data[1][48] , \cache_data[1][47] ,
         \cache_data[1][46] , \cache_data[1][45] , \cache_data[1][44] ,
         \cache_data[1][43] , \cache_data[1][42] , \cache_data[1][41] ,
         \cache_data[1][40] , \cache_data[1][39] , \cache_data[1][38] ,
         \cache_data[1][37] , \cache_data[1][36] , \cache_data[1][35] ,
         \cache_data[1][34] , \cache_data[1][33] , \cache_data[1][32] ,
         \cache_data[1][31] , \cache_data[1][30] , \cache_data[1][29] ,
         \cache_data[1][28] , \cache_data[1][27] , \cache_data[1][26] ,
         \cache_data[1][25] , \cache_data[1][24] , \cache_data[1][23] ,
         \cache_data[1][22] , \cache_data[1][21] , \cache_data[1][20] ,
         \cache_data[1][19] , \cache_data[1][18] , \cache_data[1][17] ,
         \cache_data[1][16] , \cache_data[1][15] , \cache_data[1][14] ,
         \cache_data[1][13] , \cache_data[1][12] , \cache_data[1][11] ,
         \cache_data[1][10] , \cache_data[1][9] , \cache_data[1][8] ,
         \cache_data[1][7] , \cache_data[1][6] , \cache_data[1][5] ,
         \cache_data[1][4] , \cache_data[1][3] , \cache_data[1][2] ,
         \cache_data[1][1] , \cache_data[1][0] , \cache_data[0][127] ,
         \cache_data[0][126] , \cache_data[0][125] , \cache_data[0][124] ,
         \cache_data[0][123] , \cache_data[0][122] , \cache_data[0][121] ,
         \cache_data[0][120] , \cache_data[0][119] , \cache_data[0][118] ,
         \cache_data[0][117] , \cache_data[0][116] , \cache_data[0][115] ,
         \cache_data[0][114] , \cache_data[0][113] , \cache_data[0][112] ,
         \cache_data[0][111] , \cache_data[0][110] , \cache_data[0][109] ,
         \cache_data[0][108] , \cache_data[0][107] , \cache_data[0][106] ,
         \cache_data[0][105] , \cache_data[0][104] , \cache_data[0][103] ,
         \cache_data[0][102] , \cache_data[0][101] , \cache_data[0][100] ,
         \cache_data[0][99] , \cache_data[0][98] , \cache_data[0][97] ,
         \cache_data[0][96] , \cache_data[0][95] , \cache_data[0][94] ,
         \cache_data[0][93] , \cache_data[0][92] , \cache_data[0][91] ,
         \cache_data[0][90] , \cache_data[0][89] , \cache_data[0][88] ,
         \cache_data[0][87] , \cache_data[0][86] , \cache_data[0][85] ,
         \cache_data[0][84] , \cache_data[0][83] , \cache_data[0][82] ,
         \cache_data[0][81] , \cache_data[0][80] , \cache_data[0][79] ,
         \cache_data[0][78] , \cache_data[0][77] , \cache_data[0][76] ,
         \cache_data[0][75] , \cache_data[0][74] , \cache_data[0][73] ,
         \cache_data[0][72] , \cache_data[0][71] , \cache_data[0][70] ,
         \cache_data[0][69] , \cache_data[0][68] , \cache_data[0][67] ,
         \cache_data[0][66] , \cache_data[0][65] , \cache_data[0][64] ,
         \cache_data[0][63] , \cache_data[0][62] , \cache_data[0][61] ,
         \cache_data[0][60] , \cache_data[0][59] , \cache_data[0][58] ,
         \cache_data[0][57] , \cache_data[0][56] , \cache_data[0][55] ,
         \cache_data[0][54] , \cache_data[0][53] , \cache_data[0][52] ,
         \cache_data[0][51] , \cache_data[0][50] , \cache_data[0][49] ,
         \cache_data[0][48] , \cache_data[0][47] , \cache_data[0][46] ,
         \cache_data[0][45] , \cache_data[0][44] , \cache_data[0][43] ,
         \cache_data[0][42] , \cache_data[0][41] , \cache_data[0][40] ,
         \cache_data[0][39] , \cache_data[0][38] , \cache_data[0][37] ,
         \cache_data[0][36] , \cache_data[0][35] , \cache_data[0][34] ,
         \cache_data[0][33] , \cache_data[0][32] , \cache_data[0][31] ,
         \cache_data[0][30] , \cache_data[0][29] , \cache_data[0][28] ,
         \cache_data[0][27] , \cache_data[0][26] , \cache_data[0][25] ,
         \cache_data[0][24] , \cache_data[0][23] , \cache_data[0][22] ,
         \cache_data[0][21] , \cache_data[0][20] , \cache_data[0][19] ,
         \cache_data[0][18] , \cache_data[0][17] , \cache_data[0][16] ,
         \cache_data[0][15] , \cache_data[0][14] , \cache_data[0][13] ,
         \cache_data[0][12] , \cache_data[0][11] , \cache_data[0][10] ,
         \cache_data[0][9] , \cache_data[0][8] , \cache_data[0][7] ,
         \cache_data[0][6] , \cache_data[0][5] , \cache_data[0][4] ,
         \cache_data[0][3] , \cache_data[0][2] , \cache_data[0][1] ,
         \cache_data[0][0] , rd_temp, N3426, N3427, N3429, N3430, N3432, N3433,
         N3435, N3436, N3438, N3439, N3441, N3442, N3444, N3445, N3447, N3448,
         N3450, N3451, N3453, N3454, N3456, N3457, N3459, N3460, N3462, N3463,
         N3465, N3466, N3468, N3469, N3471, N3472, N3474, N3475, N3477, N3478,
         N3480, N3481, N3483, N3484, N3486, N3487, N3489, N3490, N3492, N3493,
         N3495, N3496, N3498, N3499, N3501, N3502, N3504, N3505, N3507, N3508,
         N3510, N3511, N3513, N3514, N3516, N3517, N3519, N3520, N3522, N3523,
         N3525, N3526, N3528, N3529, N3531, N3532, N3534, N3535, N3537, N3538,
         N3540, N3541, N3543, N3544, N3546, N3547, N3549, N3550, N3552, N3553,
         N3555, N3556, N3558, N3559, N3561, N3562, N3564, N3565, N3567, N3568,
         N3570, N3571, N3573, N3574, N3576, N3577, N3579, N3580, N3582, N3583,
         N3585, N3586, N3588, N3589, N3591, N3592, N3594, N3595, N3597, N3598,
         N3600, N3601, N3603, N3604, N3606, N3607, N3609, N3610, N3612, N3613,
         N3615, N3616, N3691, N3698, n1, n3, n5, n7, n9, n11, n13, n15, n17,
         n19, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45,
         n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73,
         n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n101,
         n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, n123,
         n125, n127, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336;
  wire   [4:0] state;
  wire   [4:0] next_state;
  wire   [3:0] mem_data_cnt;
  wire   [31:0] iCache_data_wr;
  wire   [15:0] cache_valid;
  wire   [15:0] cache_dirty;
  assign addr_mem[0] = 1'b0;
  assign addr_mem[1] = 1'b0;

  drsp_1 mem_done_reg ( .ip(N3698), .ck(clk), .rb(1'b1), .s(n12324), .q(
        mem_done) );
  drsp_1 \addr_resp_tri_enable_reg[0]  ( .ip(n7408), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3616) );
  drsp_1 \addr_resp_tri_enable_reg[1]  ( .ip(n7406), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3613) );
  drsp_1 \addr_resp_tri_enable_reg[2]  ( .ip(n7404), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3610) );
  drsp_1 \addr_resp_tri_enable_reg[3]  ( .ip(n7402), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3607) );
  drsp_1 \addr_resp_tri_enable_reg[4]  ( .ip(n7400), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3604) );
  drsp_1 \addr_resp_tri_enable_reg[5]  ( .ip(n7398), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3601) );
  drsp_1 \addr_resp_tri_enable_reg[6]  ( .ip(n7396), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3598) );
  drsp_1 \addr_resp_tri_enable_reg[7]  ( .ip(n7394), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3595) );
  drsp_1 \addr_resp_tri_enable_reg[8]  ( .ip(n7376), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3592) );
  drsp_1 \addr_resp_tri_enable_reg[9]  ( .ip(n7358), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3589) );
  drsp_1 \addr_resp_tri_enable_reg[10]  ( .ip(n7340), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3586) );
  drsp_1 \addr_resp_tri_enable_reg[11]  ( .ip(n7322), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3583) );
  drsp_1 \addr_resp_tri_enable_reg[12]  ( .ip(n7304), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3580) );
  drsp_1 \addr_resp_tri_enable_reg[13]  ( .ip(n7286), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3577) );
  drsp_1 \addr_resp_tri_enable_reg[14]  ( .ip(n7268), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3574) );
  drsp_1 \addr_resp_tri_enable_reg[15]  ( .ip(n7250), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3571) );
  drsp_1 \addr_resp_tri_enable_reg[16]  ( .ip(n7232), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3568) );
  drsp_1 \addr_resp_tri_enable_reg[17]  ( .ip(n7214), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3565) );
  drsp_1 \addr_resp_tri_enable_reg[18]  ( .ip(n7196), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3562) );
  drsp_1 \addr_resp_tri_enable_reg[19]  ( .ip(n7178), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3559) );
  drsp_1 \addr_resp_tri_enable_reg[20]  ( .ip(n7160), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3556) );
  drsp_1 \addr_resp_tri_enable_reg[21]  ( .ip(n7142), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3553) );
  drsp_1 \addr_resp_tri_enable_reg[22]  ( .ip(n7124), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3550) );
  drsp_1 \addr_resp_tri_enable_reg[23]  ( .ip(n7106), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3547) );
  drsp_1 \addr_resp_tri_enable_reg[24]  ( .ip(n7088), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3544) );
  drsp_1 \addr_resp_tri_enable_reg[25]  ( .ip(n7070), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3541) );
  drsp_1 \addr_resp_tri_enable_reg[26]  ( .ip(n7052), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3538) );
  drsp_1 \addr_resp_tri_enable_reg[27]  ( .ip(n7034), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3535) );
  drsp_1 \addr_resp_tri_enable_reg[28]  ( .ip(n7016), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3532) );
  drsp_1 \addr_resp_tri_enable_reg[29]  ( .ip(n6998), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3529) );
  drsp_1 \addr_resp_tri_enable_reg[30]  ( .ip(n6980), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3526) );
  drsp_1 \addr_resp_tri_enable_reg[31]  ( .ip(n6962), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3523) );
  drsp_1 rd_temp_reg ( .ip(n6945), .ck(clk), .rb(1'b1), .s(n12336), .q(rd_temp) );
  drsp_1 \state_reg[0]  ( .ip(next_state[0]), .ck(clk), .rb(1'b1), .s(n12335), 
        .q(state[0]) );
  drsp_1 busy_reg ( .ip(N3691), .ck(clk), .rb(1'b1), .s(n12335), .q(busy) );
  drsp_1 \data_rd_tri_enable_reg[0]  ( .ip(n6943), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3520) );
  drsp_1 \data_rd_tri_enable_reg[1]  ( .ip(n6941), .ck(clk), .rb(1'b1), .s(rst), .q(N3517) );
  drsp_1 \data_rd_tri_enable_reg[2]  ( .ip(n6939), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3514) );
  drsp_1 \data_rd_tri_enable_reg[3]  ( .ip(n6937), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3511) );
  drsp_1 \data_rd_tri_enable_reg[4]  ( .ip(n6935), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3508) );
  drsp_1 \data_rd_tri_enable_reg[5]  ( .ip(n6933), .ck(clk), .rb(1'b1), .s(rst), .q(N3505) );
  drsp_1 \data_rd_tri_enable_reg[6]  ( .ip(n6931), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3502) );
  drsp_1 \data_rd_tri_enable_reg[7]  ( .ip(n6929), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3499) );
  drsp_1 \data_rd_tri_enable_reg[8]  ( .ip(n6927), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3496) );
  drsp_1 \data_rd_tri_enable_reg[9]  ( .ip(n6925), .ck(clk), .rb(1'b1), .s(rst), .q(N3493) );
  drsp_1 \data_rd_tri_enable_reg[10]  ( .ip(n6923), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3490) );
  drsp_1 \data_rd_tri_enable_reg[11]  ( .ip(n6921), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3487) );
  drsp_1 \data_rd_tri_enable_reg[12]  ( .ip(n6919), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3484) );
  drsp_1 \data_rd_tri_enable_reg[13]  ( .ip(n6917), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3481) );
  drsp_1 \data_rd_tri_enable_reg[14]  ( .ip(n6915), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3478) );
  drsp_1 \data_rd_tri_enable_reg[15]  ( .ip(n6913), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3475) );
  drsp_1 \data_rd_tri_enable_reg[16]  ( .ip(n6911), .ck(clk), .rb(1'b1), .s(
        n12324), .q(N3472) );
  drsp_1 \data_rd_tri_enable_reg[17]  ( .ip(n6909), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3469) );
  drsp_1 \data_rd_tri_enable_reg[18]  ( .ip(n6907), .ck(clk), .rb(1'b1), .s(
        rst), .q(N3466) );
  drsp_1 \data_rd_tri_enable_reg[19]  ( .ip(n6905), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3463) );
  drsp_1 \data_rd_tri_enable_reg[20]  ( .ip(n6903), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3460) );
  drsp_1 \data_rd_tri_enable_reg[21]  ( .ip(n6901), .ck(clk), .rb(1'b1), .s(
        n12334), .q(N3457) );
  drsp_1 \data_rd_tri_enable_reg[22]  ( .ip(n6899), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3454) );
  drsp_1 \data_rd_tri_enable_reg[23]  ( .ip(n6897), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3451) );
  drsp_1 \data_rd_tri_enable_reg[24]  ( .ip(n6895), .ck(clk), .rb(1'b1), .s(
        n12335), .q(N3448) );
  drsp_1 \data_rd_tri_enable_reg[25]  ( .ip(n6893), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3445) );
  drsp_1 \data_rd_tri_enable_reg[26]  ( .ip(n6891), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3442) );
  drsp_1 \data_rd_tri_enable_reg[27]  ( .ip(n6889), .ck(clk), .rb(1'b1), .s(
        n12336), .q(N3439) );
  drsp_1 \data_rd_tri_enable_reg[28]  ( .ip(n6887), .ck(clk), .rb(1'b1), .s(
        n12324), .q(N3436) );
  drsp_1 \data_rd_tri_enable_reg[29]  ( .ip(n6885), .ck(clk), .rb(1'b1), .s(
        n12324), .q(N3433) );
  drsp_1 \data_rd_tri_enable_reg[30]  ( .ip(n6883), .ck(clk), .rb(1'b1), .s(
        n12324), .q(N3430) );
  drsp_1 \data_rd_tri_enable_reg[31]  ( .ip(n6881), .ck(clk), .rb(1'b1), .s(
        n12324), .q(N3427) );
  drp_1 \state_reg[4]  ( .ip(n12323), .ck(clk), .rb(n12326), .q(state[4]) );
  drp_1 miss_reg ( .ip(n7412), .ck(clk), .rb(n12326), .q(miss) );
  drp_1 valid_reg ( .ip(n7411), .ck(clk), .rb(n12326), .q(valid) );
  drp_1 dirty_reg ( .ip(n7410), .ck(clk), .rb(n12326), .q(dirty) );
  drp_1 hit_reg ( .ip(n6864), .ck(clk), .rb(n12326), .q(hit) );
  drp_1 \state_reg[3]  ( .ip(n12325), .ck(clk), .rb(n12326), .q(state[3]) );
  drp_1 \state_reg[2]  ( .ip(next_state[2]), .ck(clk), .rb(n12326), .q(
        state[2]) );
  drp_1 \state_reg[1]  ( .ip(next_state[1]), .ck(clk), .rb(n12333), .q(
        state[1]) );
  drp_1 \mem_data_cnt_reg[2]  ( .ip(n7415), .ck(clk), .rb(n12333), .q(
        mem_data_cnt[2]) );
  drp_1 \mem_data_cnt_reg[3]  ( .ip(n7416), .ck(clk), .rb(n12333), .q(
        mem_data_cnt[3]) );
  drp_1 \cache_valid_reg[0]  ( .ip(n7393), .ck(clk), .rb(n12333), .q(
        cache_valid[0]) );
  drp_1 \cache_valid_reg[1]  ( .ip(n7392), .ck(clk), .rb(n12333), .q(
        cache_valid[1]) );
  drp_1 \cache_valid_reg[2]  ( .ip(n7391), .ck(clk), .rb(n12333), .q(
        cache_valid[2]) );
  drp_1 \cache_valid_reg[3]  ( .ip(n7390), .ck(clk), .rb(n12333), .q(
        cache_valid[3]) );
  drp_1 \cache_valid_reg[4]  ( .ip(n7389), .ck(clk), .rb(n12333), .q(
        cache_valid[4]) );
  drp_1 \cache_valid_reg[5]  ( .ip(n7388), .ck(clk), .rb(n12333), .q(
        cache_valid[5]) );
  drp_1 \cache_valid_reg[6]  ( .ip(n7387), .ck(clk), .rb(n12333), .q(
        cache_valid[6]) );
  drp_1 \cache_valid_reg[7]  ( .ip(n7386), .ck(clk), .rb(n12333), .q(
        cache_valid[7]) );
  drp_1 \cache_valid_reg[8]  ( .ip(n7385), .ck(clk), .rb(n12333), .q(
        cache_valid[8]) );
  drp_1 \cache_valid_reg[9]  ( .ip(n7384), .ck(clk), .rb(n12327), .q(
        cache_valid[9]) );
  drp_1 \cache_valid_reg[10]  ( .ip(n7383), .ck(clk), .rb(n12328), .q(
        cache_valid[10]) );
  drp_1 \cache_valid_reg[11]  ( .ip(n7382), .ck(clk), .rb(n12329), .q(
        cache_valid[11]) );
  drp_1 \cache_valid_reg[12]  ( .ip(n7381), .ck(clk), .rb(n12330), .q(
        cache_valid[12]) );
  drp_1 \cache_valid_reg[13]  ( .ip(n7380), .ck(clk), .rb(n12331), .q(
        cache_valid[13]) );
  drp_1 \cache_valid_reg[14]  ( .ip(n7379), .ck(clk), .rb(n12332), .q(
        cache_valid[14]) );
  drp_1 \cache_valid_reg[15]  ( .ip(n7378), .ck(clk), .rb(n12332), .q(
        cache_valid[15]) );
  drp_1 rdy_reg ( .ip(n12323), .ck(clk), .rb(n12327), .q(rdy) );
  drp_1 \cache_dirty_reg[0]  ( .ip(n6880), .ck(clk), .rb(n12328), .q(
        cache_dirty[0]) );
  drp_1 \cache_dirty_reg[1]  ( .ip(n6879), .ck(clk), .rb(n12329), .q(
        cache_dirty[1]) );
  drp_1 \cache_dirty_reg[2]  ( .ip(n6878), .ck(clk), .rb(n12330), .q(
        cache_dirty[2]) );
  drp_1 \cache_dirty_reg[3]  ( .ip(n6877), .ck(clk), .rb(n12331), .q(
        cache_dirty[3]) );
  drp_1 \cache_dirty_reg[4]  ( .ip(n6876), .ck(clk), .rb(n12330), .q(
        cache_dirty[4]) );
  drp_1 \cache_dirty_reg[5]  ( .ip(n6875), .ck(clk), .rb(n12331), .q(
        cache_dirty[5]) );
  drp_1 \cache_dirty_reg[6]  ( .ip(n6874), .ck(clk), .rb(n12332), .q(
        cache_dirty[6]) );
  drp_1 \cache_dirty_reg[7]  ( .ip(n6873), .ck(clk), .rb(n12327), .q(
        cache_dirty[7]) );
  drp_1 \cache_dirty_reg[8]  ( .ip(n6872), .ck(clk), .rb(n12328), .q(
        cache_dirty[8]) );
  drp_1 \cache_dirty_reg[9]  ( .ip(n6871), .ck(clk), .rb(n12329), .q(
        cache_dirty[9]) );
  drp_1 \cache_dirty_reg[10]  ( .ip(n6870), .ck(clk), .rb(n12330), .q(
        cache_dirty[10]) );
  drp_1 \cache_dirty_reg[11]  ( .ip(n6869), .ck(clk), .rb(n12331), .q(
        cache_dirty[11]) );
  drp_1 \cache_dirty_reg[12]  ( .ip(n6868), .ck(clk), .rb(n12332), .q(
        cache_dirty[12]) );
  drp_1 \cache_dirty_reg[13]  ( .ip(n6867), .ck(clk), .rb(n12327), .q(
        cache_dirty[13]) );
  drp_1 \cache_dirty_reg[14]  ( .ip(n6866), .ck(clk), .rb(n12328), .q(
        cache_dirty[14]) );
  drp_1 \cache_dirty_reg[15]  ( .ip(n6865), .ck(clk), .rb(n12329), .q(
        cache_dirty[15]) );
  drp_1 \addr_mem_reg[2]  ( .ip(n4781), .ck(clk), .rb(n12332), .q(addr_mem[2])
         );
  drp_1 \addr_mem_reg[3]  ( .ip(n4780), .ck(clk), .rb(n12332), .q(addr_mem[3])
         );
  drp_1 \addr_mem_reg[4]  ( .ip(n4779), .ck(clk), .rb(n12332), .q(addr_mem[4])
         );
  drp_1 \addr_mem_reg[5]  ( .ip(n4778), .ck(clk), .rb(n12332), .q(addr_mem[5])
         );
  drp_1 \addr_mem_reg[6]  ( .ip(n4777), .ck(clk), .rb(n12332), .q(addr_mem[6])
         );
  drp_1 \addr_mem_reg[7]  ( .ip(n4776), .ck(clk), .rb(n12332), .q(addr_mem[7])
         );
  drp_1 wr_mem_reg ( .ip(n7414), .ck(clk), .rb(n12332), .q(wr_mem) );
  drp_1 rd_mem_reg ( .ip(n7413), .ck(clk), .rb(n12332), .q(rd_mem) );
  drp_1 \addr_mem_reg[8]  ( .ip(n4775), .ck(clk), .rb(n12332), .q(addr_mem[8])
         );
  drp_1 \addr_mem_reg[9]  ( .ip(n4774), .ck(clk), .rb(n12332), .q(addr_mem[9])
         );
  drp_1 \addr_mem_reg[10]  ( .ip(n4773), .ck(clk), .rb(n12332), .q(
        addr_mem[10]) );
  drp_1 \addr_mem_reg[11]  ( .ip(n4772), .ck(clk), .rb(n12332), .q(
        addr_mem[11]) );
  drp_1 \addr_mem_reg[12]  ( .ip(n4771), .ck(clk), .rb(n12331), .q(
        addr_mem[12]) );
  drp_1 \addr_mem_reg[13]  ( .ip(n4770), .ck(clk), .rb(n12331), .q(
        addr_mem[13]) );
  drp_1 \addr_mem_reg[14]  ( .ip(n4769), .ck(clk), .rb(n12331), .q(
        addr_mem[14]) );
  drp_1 \addr_mem_reg[15]  ( .ip(n4768), .ck(clk), .rb(n12331), .q(
        addr_mem[15]) );
  drp_1 \addr_mem_reg[16]  ( .ip(n4767), .ck(clk), .rb(n12331), .q(
        addr_mem[16]) );
  drp_1 \addr_mem_reg[17]  ( .ip(n4766), .ck(clk), .rb(n12331), .q(
        addr_mem[17]) );
  drp_1 \addr_mem_reg[18]  ( .ip(n4765), .ck(clk), .rb(n12331), .q(
        addr_mem[18]) );
  drp_1 \addr_mem_reg[19]  ( .ip(n4764), .ck(clk), .rb(n12331), .q(
        addr_mem[19]) );
  drp_1 \addr_mem_reg[20]  ( .ip(n4763), .ck(clk), .rb(n12331), .q(
        addr_mem[20]) );
  drp_1 \addr_mem_reg[21]  ( .ip(n4762), .ck(clk), .rb(n12331), .q(
        addr_mem[21]) );
  drp_1 \addr_mem_reg[22]  ( .ip(n4761), .ck(clk), .rb(n12331), .q(
        addr_mem[22]) );
  drp_1 \addr_mem_reg[23]  ( .ip(n4760), .ck(clk), .rb(n12331), .q(
        addr_mem[23]) );
  drp_1 \addr_mem_reg[24]  ( .ip(n4759), .ck(clk), .rb(n12330), .q(
        addr_mem[24]) );
  drp_1 \addr_mem_reg[25]  ( .ip(n4758), .ck(clk), .rb(n12330), .q(
        addr_mem[25]) );
  drp_1 \addr_mem_reg[26]  ( .ip(n4757), .ck(clk), .rb(n12330), .q(
        addr_mem[26]) );
  drp_1 \addr_mem_reg[27]  ( .ip(n4756), .ck(clk), .rb(n12330), .q(
        addr_mem[27]) );
  drp_1 \addr_mem_reg[28]  ( .ip(n4755), .ck(clk), .rb(n12330), .q(
        addr_mem[28]) );
  drp_1 \addr_mem_reg[29]  ( .ip(n4754), .ck(clk), .rb(n12330), .q(
        addr_mem[29]) );
  drp_1 \addr_mem_reg[30]  ( .ip(n4753), .ck(clk), .rb(n12330), .q(
        addr_mem[30]) );
  drp_1 \addr_mem_reg[31]  ( .ip(n4752), .ck(clk), .rb(n12330), .q(
        addr_mem[31]) );
  dp_1 \addr_resp_reg[0]  ( .ip(n7409), .ck(clk), .q(N3615) );
  dp_1 \addr_resp_reg[1]  ( .ip(n7407), .ck(clk), .q(N3612) );
  dp_1 \addr_resp_reg[2]  ( .ip(n7405), .ck(clk), .q(N3609) );
  dp_1 \addr_resp_reg[3]  ( .ip(n7403), .ck(clk), .q(N3606) );
  dp_1 \addr_resp_reg[4]  ( .ip(n7401), .ck(clk), .q(N3603) );
  dp_1 \addr_resp_reg[5]  ( .ip(n7399), .ck(clk), .q(N3600) );
  dp_1 \addr_resp_reg[6]  ( .ip(n7397), .ck(clk), .q(N3597) );
  dp_1 \addr_resp_reg[7]  ( .ip(n7395), .ck(clk), .q(N3594) );
  dp_1 \addr_resp_reg[8]  ( .ip(n7377), .ck(clk), .q(N3591) );
  dp_1 \addr_resp_reg[9]  ( .ip(n7359), .ck(clk), .q(N3588) );
  dp_1 \addr_resp_reg[10]  ( .ip(n7341), .ck(clk), .q(N3585) );
  dp_1 \addr_resp_reg[11]  ( .ip(n7323), .ck(clk), .q(N3582) );
  dp_1 \addr_resp_reg[12]  ( .ip(n7305), .ck(clk), .q(N3579) );
  dp_1 \addr_resp_reg[13]  ( .ip(n7287), .ck(clk), .q(N3576) );
  dp_1 \addr_resp_reg[14]  ( .ip(n7269), .ck(clk), .q(N3573) );
  dp_1 \addr_resp_reg[15]  ( .ip(n7251), .ck(clk), .q(N3570) );
  dp_1 \addr_resp_reg[16]  ( .ip(n7233), .ck(clk), .q(N3567) );
  dp_1 \addr_resp_reg[17]  ( .ip(n7215), .ck(clk), .q(N3564) );
  dp_1 \addr_resp_reg[18]  ( .ip(n7197), .ck(clk), .q(N3561) );
  dp_1 \addr_resp_reg[19]  ( .ip(n7179), .ck(clk), .q(N3558) );
  dp_1 \addr_resp_reg[20]  ( .ip(n7161), .ck(clk), .q(N3555) );
  dp_1 \addr_resp_reg[21]  ( .ip(n7143), .ck(clk), .q(N3552) );
  dp_1 \addr_resp_reg[22]  ( .ip(n7125), .ck(clk), .q(N3549) );
  dp_1 \addr_resp_reg[23]  ( .ip(n7107), .ck(clk), .q(N3546) );
  dp_1 \addr_resp_reg[24]  ( .ip(n7089), .ck(clk), .q(N3543) );
  dp_1 \addr_resp_reg[25]  ( .ip(n7071), .ck(clk), .q(N3540) );
  dp_1 \addr_resp_reg[26]  ( .ip(n7053), .ck(clk), .q(N3537) );
  dp_1 \addr_resp_reg[27]  ( .ip(n7035), .ck(clk), .q(N3534) );
  dp_1 \addr_resp_reg[28]  ( .ip(n7017), .ck(clk), .q(N3531) );
  dp_1 \addr_resp_reg[29]  ( .ip(n6999), .ck(clk), .q(N3528) );
  dp_1 \addr_resp_reg[30]  ( .ip(n6981), .ck(clk), .q(N3525) );
  dp_1 \addr_resp_reg[31]  ( .ip(n6963), .ck(clk), .q(N3522) );
  dp_1 \data_wr_mem_reg[0]  ( .ip(n7448), .ck(clk), .q(data_wr_mem[0]) );
  dp_1 \data_wr_mem_reg[1]  ( .ip(n7447), .ck(clk), .q(data_wr_mem[1]) );
  dp_1 \data_wr_mem_reg[2]  ( .ip(n7446), .ck(clk), .q(data_wr_mem[2]) );
  dp_1 \data_wr_mem_reg[3]  ( .ip(n7445), .ck(clk), .q(data_wr_mem[3]) );
  dp_1 \data_wr_mem_reg[4]  ( .ip(n7444), .ck(clk), .q(data_wr_mem[4]) );
  dp_1 \data_wr_mem_reg[5]  ( .ip(n7443), .ck(clk), .q(data_wr_mem[5]) );
  dp_1 \data_wr_mem_reg[6]  ( .ip(n7442), .ck(clk), .q(data_wr_mem[6]) );
  dp_1 \data_wr_mem_reg[7]  ( .ip(n7441), .ck(clk), .q(data_wr_mem[7]) );
  dp_1 \data_wr_mem_reg[8]  ( .ip(n7440), .ck(clk), .q(data_wr_mem[8]) );
  dp_1 \data_wr_mem_reg[9]  ( .ip(n7439), .ck(clk), .q(data_wr_mem[9]) );
  dp_1 \data_wr_mem_reg[10]  ( .ip(n7438), .ck(clk), .q(data_wr_mem[10]) );
  dp_1 \data_wr_mem_reg[11]  ( .ip(n7437), .ck(clk), .q(data_wr_mem[11]) );
  dp_1 \data_wr_mem_reg[12]  ( .ip(n7436), .ck(clk), .q(data_wr_mem[12]) );
  dp_1 \data_wr_mem_reg[13]  ( .ip(n7435), .ck(clk), .q(data_wr_mem[13]) );
  dp_1 \data_wr_mem_reg[14]  ( .ip(n7434), .ck(clk), .q(data_wr_mem[14]) );
  dp_1 \data_wr_mem_reg[15]  ( .ip(n7433), .ck(clk), .q(data_wr_mem[15]) );
  dp_1 \data_wr_mem_reg[16]  ( .ip(n7432), .ck(clk), .q(data_wr_mem[16]) );
  dp_1 \data_wr_mem_reg[17]  ( .ip(n7431), .ck(clk), .q(data_wr_mem[17]) );
  dp_1 \data_wr_mem_reg[18]  ( .ip(n7430), .ck(clk), .q(data_wr_mem[18]) );
  dp_1 \data_wr_mem_reg[19]  ( .ip(n7429), .ck(clk), .q(data_wr_mem[19]) );
  dp_1 \data_wr_mem_reg[20]  ( .ip(n7428), .ck(clk), .q(data_wr_mem[20]) );
  dp_1 \data_wr_mem_reg[21]  ( .ip(n7427), .ck(clk), .q(data_wr_mem[21]) );
  dp_1 \data_wr_mem_reg[22]  ( .ip(n7426), .ck(clk), .q(data_wr_mem[22]) );
  dp_1 \data_wr_mem_reg[23]  ( .ip(n7425), .ck(clk), .q(data_wr_mem[23]) );
  dp_1 \data_wr_mem_reg[24]  ( .ip(n7424), .ck(clk), .q(data_wr_mem[24]) );
  dp_1 \data_wr_mem_reg[25]  ( .ip(n7423), .ck(clk), .q(data_wr_mem[25]) );
  dp_1 \data_wr_mem_reg[26]  ( .ip(n7422), .ck(clk), .q(data_wr_mem[26]) );
  dp_1 \data_wr_mem_reg[27]  ( .ip(n7421), .ck(clk), .q(data_wr_mem[27]) );
  dp_1 \data_wr_mem_reg[28]  ( .ip(n7420), .ck(clk), .q(data_wr_mem[28]) );
  dp_1 \data_wr_mem_reg[29]  ( .ip(n7419), .ck(clk), .q(data_wr_mem[29]) );
  dp_1 \data_wr_mem_reg[30]  ( .ip(n7418), .ck(clk), .q(data_wr_mem[30]) );
  dp_1 \data_wr_mem_reg[31]  ( .ip(n7417), .ck(clk), .q(data_wr_mem[31]) );
  dp_1 \cache_tag_reg[0][0]  ( .ip(n7375), .ck(clk), .q(\cache_tag[0][0] ) );
  dp_1 \cache_tag_reg[0][1]  ( .ip(n7357), .ck(clk), .q(\cache_tag[0][1] ) );
  dp_1 \cache_tag_reg[0][2]  ( .ip(n7339), .ck(clk), .q(\cache_tag[0][2] ) );
  dp_1 \cache_tag_reg[0][3]  ( .ip(n7321), .ck(clk), .q(\cache_tag[0][3] ) );
  dp_1 \cache_tag_reg[0][4]  ( .ip(n7303), .ck(clk), .q(\cache_tag[0][4] ) );
  dp_1 \cache_tag_reg[0][5]  ( .ip(n7285), .ck(clk), .q(\cache_tag[0][5] ) );
  dp_1 \cache_tag_reg[0][6]  ( .ip(n7267), .ck(clk), .q(\cache_tag[0][6] ) );
  dp_1 \cache_tag_reg[0][7]  ( .ip(n7249), .ck(clk), .q(\cache_tag[0][7] ) );
  dp_1 \cache_tag_reg[0][8]  ( .ip(n7231), .ck(clk), .q(\cache_tag[0][8] ) );
  dp_1 \cache_tag_reg[0][9]  ( .ip(n7213), .ck(clk), .q(\cache_tag[0][9] ) );
  dp_1 \cache_tag_reg[0][10]  ( .ip(n7195), .ck(clk), .q(\cache_tag[0][10] )
         );
  dp_1 \cache_tag_reg[0][11]  ( .ip(n7177), .ck(clk), .q(\cache_tag[0][11] )
         );
  dp_1 \cache_tag_reg[0][12]  ( .ip(n7159), .ck(clk), .q(\cache_tag[0][12] )
         );
  dp_1 \cache_tag_reg[0][13]  ( .ip(n7141), .ck(clk), .q(\cache_tag[0][13] )
         );
  dp_1 \cache_tag_reg[0][14]  ( .ip(n7123), .ck(clk), .q(\cache_tag[0][14] )
         );
  dp_1 \cache_tag_reg[0][15]  ( .ip(n7105), .ck(clk), .q(\cache_tag[0][15] )
         );
  dp_1 \cache_tag_reg[0][16]  ( .ip(n7087), .ck(clk), .q(\cache_tag[0][16] )
         );
  dp_1 \cache_tag_reg[0][17]  ( .ip(n7069), .ck(clk), .q(\cache_tag[0][17] )
         );
  dp_1 \cache_tag_reg[0][18]  ( .ip(n7051), .ck(clk), .q(\cache_tag[0][18] )
         );
  dp_1 \cache_tag_reg[0][19]  ( .ip(n7033), .ck(clk), .q(\cache_tag[0][19] )
         );
  dp_1 \cache_tag_reg[0][20]  ( .ip(n7015), .ck(clk), .q(\cache_tag[0][20] )
         );
  dp_1 \cache_tag_reg[0][21]  ( .ip(n6997), .ck(clk), .q(\cache_tag[0][21] )
         );
  dp_1 \cache_tag_reg[0][22]  ( .ip(n6979), .ck(clk), .q(\cache_tag[0][22] )
         );
  dp_1 \cache_tag_reg[0][23]  ( .ip(n6961), .ck(clk), .q(\cache_tag[0][23] )
         );
  dp_1 \cache_tag_reg[1][0]  ( .ip(n7374), .ck(clk), .q(\cache_tag[1][0] ) );
  dp_1 \cache_tag_reg[1][1]  ( .ip(n7356), .ck(clk), .q(\cache_tag[1][1] ) );
  dp_1 \cache_tag_reg[1][2]  ( .ip(n7338), .ck(clk), .q(\cache_tag[1][2] ) );
  dp_1 \cache_tag_reg[1][3]  ( .ip(n7320), .ck(clk), .q(\cache_tag[1][3] ) );
  dp_1 \cache_tag_reg[1][4]  ( .ip(n7302), .ck(clk), .q(\cache_tag[1][4] ) );
  dp_1 \cache_tag_reg[1][5]  ( .ip(n7284), .ck(clk), .q(\cache_tag[1][5] ) );
  dp_1 \cache_tag_reg[1][6]  ( .ip(n7266), .ck(clk), .q(\cache_tag[1][6] ) );
  dp_1 \cache_tag_reg[1][7]  ( .ip(n7248), .ck(clk), .q(\cache_tag[1][7] ) );
  dp_1 \cache_tag_reg[1][8]  ( .ip(n7230), .ck(clk), .q(\cache_tag[1][8] ) );
  dp_1 \cache_tag_reg[1][9]  ( .ip(n7212), .ck(clk), .q(\cache_tag[1][9] ) );
  dp_1 \cache_tag_reg[1][10]  ( .ip(n7194), .ck(clk), .q(\cache_tag[1][10] )
         );
  dp_1 \cache_tag_reg[1][11]  ( .ip(n7176), .ck(clk), .q(\cache_tag[1][11] )
         );
  dp_1 \cache_tag_reg[1][12]  ( .ip(n7158), .ck(clk), .q(\cache_tag[1][12] )
         );
  dp_1 \cache_tag_reg[1][13]  ( .ip(n7140), .ck(clk), .q(\cache_tag[1][13] )
         );
  dp_1 \cache_tag_reg[1][14]  ( .ip(n7122), .ck(clk), .q(\cache_tag[1][14] )
         );
  dp_1 \cache_tag_reg[1][15]  ( .ip(n7104), .ck(clk), .q(\cache_tag[1][15] )
         );
  dp_1 \cache_tag_reg[1][16]  ( .ip(n7086), .ck(clk), .q(\cache_tag[1][16] )
         );
  dp_1 \cache_tag_reg[1][17]  ( .ip(n7068), .ck(clk), .q(\cache_tag[1][17] )
         );
  dp_1 \cache_tag_reg[1][18]  ( .ip(n7050), .ck(clk), .q(\cache_tag[1][18] )
         );
  dp_1 \cache_tag_reg[1][19]  ( .ip(n7032), .ck(clk), .q(\cache_tag[1][19] )
         );
  dp_1 \cache_tag_reg[1][20]  ( .ip(n7014), .ck(clk), .q(\cache_tag[1][20] )
         );
  dp_1 \cache_tag_reg[1][21]  ( .ip(n6996), .ck(clk), .q(\cache_tag[1][21] )
         );
  dp_1 \cache_tag_reg[1][22]  ( .ip(n6978), .ck(clk), .q(\cache_tag[1][22] )
         );
  dp_1 \cache_tag_reg[1][23]  ( .ip(n6960), .ck(clk), .q(\cache_tag[1][23] )
         );
  dp_1 \cache_tag_reg[2][0]  ( .ip(n7373), .ck(clk), .q(\cache_tag[2][0] ) );
  dp_1 \cache_tag_reg[2][1]  ( .ip(n7355), .ck(clk), .q(\cache_tag[2][1] ) );
  dp_1 \cache_tag_reg[2][2]  ( .ip(n7337), .ck(clk), .q(\cache_tag[2][2] ) );
  dp_1 \cache_tag_reg[2][3]  ( .ip(n7319), .ck(clk), .q(\cache_tag[2][3] ) );
  dp_1 \cache_tag_reg[2][4]  ( .ip(n7301), .ck(clk), .q(\cache_tag[2][4] ) );
  dp_1 \cache_tag_reg[2][5]  ( .ip(n7283), .ck(clk), .q(\cache_tag[2][5] ) );
  dp_1 \cache_tag_reg[2][6]  ( .ip(n7265), .ck(clk), .q(\cache_tag[2][6] ) );
  dp_1 \cache_tag_reg[2][7]  ( .ip(n7247), .ck(clk), .q(\cache_tag[2][7] ) );
  dp_1 \cache_tag_reg[2][8]  ( .ip(n7229), .ck(clk), .q(\cache_tag[2][8] ) );
  dp_1 \cache_tag_reg[2][9]  ( .ip(n7211), .ck(clk), .q(\cache_tag[2][9] ) );
  dp_1 \cache_tag_reg[2][10]  ( .ip(n7193), .ck(clk), .q(\cache_tag[2][10] )
         );
  dp_1 \cache_tag_reg[2][11]  ( .ip(n7175), .ck(clk), .q(\cache_tag[2][11] )
         );
  dp_1 \cache_tag_reg[2][12]  ( .ip(n7157), .ck(clk), .q(\cache_tag[2][12] )
         );
  dp_1 \cache_tag_reg[2][13]  ( .ip(n7139), .ck(clk), .q(\cache_tag[2][13] )
         );
  dp_1 \cache_tag_reg[2][14]  ( .ip(n7121), .ck(clk), .q(\cache_tag[2][14] )
         );
  dp_1 \cache_tag_reg[2][15]  ( .ip(n7103), .ck(clk), .q(\cache_tag[2][15] )
         );
  dp_1 \cache_tag_reg[2][16]  ( .ip(n7085), .ck(clk), .q(\cache_tag[2][16] )
         );
  dp_1 \cache_tag_reg[2][17]  ( .ip(n7067), .ck(clk), .q(\cache_tag[2][17] )
         );
  dp_1 \cache_tag_reg[2][18]  ( .ip(n7049), .ck(clk), .q(\cache_tag[2][18] )
         );
  dp_1 \cache_tag_reg[2][19]  ( .ip(n7031), .ck(clk), .q(\cache_tag[2][19] )
         );
  dp_1 \cache_tag_reg[2][20]  ( .ip(n7013), .ck(clk), .q(\cache_tag[2][20] )
         );
  dp_1 \cache_tag_reg[2][21]  ( .ip(n6995), .ck(clk), .q(\cache_tag[2][21] )
         );
  dp_1 \cache_tag_reg[2][22]  ( .ip(n6977), .ck(clk), .q(\cache_tag[2][22] )
         );
  dp_1 \cache_tag_reg[2][23]  ( .ip(n6959), .ck(clk), .q(\cache_tag[2][23] )
         );
  dp_1 \cache_tag_reg[3][0]  ( .ip(n7372), .ck(clk), .q(\cache_tag[3][0] ) );
  dp_1 \cache_tag_reg[3][1]  ( .ip(n7354), .ck(clk), .q(\cache_tag[3][1] ) );
  dp_1 \cache_tag_reg[3][2]  ( .ip(n7336), .ck(clk), .q(\cache_tag[3][2] ) );
  dp_1 \cache_tag_reg[3][3]  ( .ip(n7318), .ck(clk), .q(\cache_tag[3][3] ) );
  dp_1 \cache_tag_reg[3][4]  ( .ip(n7300), .ck(clk), .q(\cache_tag[3][4] ) );
  dp_1 \cache_tag_reg[3][5]  ( .ip(n7282), .ck(clk), .q(\cache_tag[3][5] ) );
  dp_1 \cache_tag_reg[3][6]  ( .ip(n7264), .ck(clk), .q(\cache_tag[3][6] ) );
  dp_1 \cache_tag_reg[3][7]  ( .ip(n7246), .ck(clk), .q(\cache_tag[3][7] ) );
  dp_1 \cache_tag_reg[3][8]  ( .ip(n7228), .ck(clk), .q(\cache_tag[3][8] ) );
  dp_1 \cache_tag_reg[3][9]  ( .ip(n7210), .ck(clk), .q(\cache_tag[3][9] ) );
  dp_1 \cache_tag_reg[3][10]  ( .ip(n7192), .ck(clk), .q(\cache_tag[3][10] )
         );
  dp_1 \cache_tag_reg[3][11]  ( .ip(n7174), .ck(clk), .q(\cache_tag[3][11] )
         );
  dp_1 \cache_tag_reg[3][12]  ( .ip(n7156), .ck(clk), .q(\cache_tag[3][12] )
         );
  dp_1 \cache_tag_reg[3][13]  ( .ip(n7138), .ck(clk), .q(\cache_tag[3][13] )
         );
  dp_1 \cache_tag_reg[3][14]  ( .ip(n7120), .ck(clk), .q(\cache_tag[3][14] )
         );
  dp_1 \cache_tag_reg[3][15]  ( .ip(n7102), .ck(clk), .q(\cache_tag[3][15] )
         );
  dp_1 \cache_tag_reg[3][16]  ( .ip(n7084), .ck(clk), .q(\cache_tag[3][16] )
         );
  dp_1 \cache_tag_reg[3][17]  ( .ip(n7066), .ck(clk), .q(\cache_tag[3][17] )
         );
  dp_1 \cache_tag_reg[3][18]  ( .ip(n7048), .ck(clk), .q(\cache_tag[3][18] )
         );
  dp_1 \cache_tag_reg[3][19]  ( .ip(n7030), .ck(clk), .q(\cache_tag[3][19] )
         );
  dp_1 \cache_tag_reg[3][20]  ( .ip(n7012), .ck(clk), .q(\cache_tag[3][20] )
         );
  dp_1 \cache_tag_reg[3][21]  ( .ip(n6994), .ck(clk), .q(\cache_tag[3][21] )
         );
  dp_1 \cache_tag_reg[3][22]  ( .ip(n6976), .ck(clk), .q(\cache_tag[3][22] )
         );
  dp_1 \cache_tag_reg[3][23]  ( .ip(n6958), .ck(clk), .q(\cache_tag[3][23] )
         );
  dp_1 \cache_tag_reg[4][0]  ( .ip(n7371), .ck(clk), .q(\cache_tag[4][0] ) );
  dp_1 \cache_tag_reg[4][1]  ( .ip(n7353), .ck(clk), .q(\cache_tag[4][1] ) );
  dp_1 \cache_tag_reg[4][2]  ( .ip(n7335), .ck(clk), .q(\cache_tag[4][2] ) );
  dp_1 \cache_tag_reg[4][3]  ( .ip(n7317), .ck(clk), .q(\cache_tag[4][3] ) );
  dp_1 \cache_tag_reg[4][4]  ( .ip(n7299), .ck(clk), .q(\cache_tag[4][4] ) );
  dp_1 \cache_tag_reg[4][5]  ( .ip(n7281), .ck(clk), .q(\cache_tag[4][5] ) );
  dp_1 \cache_tag_reg[4][6]  ( .ip(n7263), .ck(clk), .q(\cache_tag[4][6] ) );
  dp_1 \cache_tag_reg[4][7]  ( .ip(n7245), .ck(clk), .q(\cache_tag[4][7] ) );
  dp_1 \cache_tag_reg[4][8]  ( .ip(n7227), .ck(clk), .q(\cache_tag[4][8] ) );
  dp_1 \cache_tag_reg[4][9]  ( .ip(n7209), .ck(clk), .q(\cache_tag[4][9] ) );
  dp_1 \cache_tag_reg[4][10]  ( .ip(n7191), .ck(clk), .q(\cache_tag[4][10] )
         );
  dp_1 \cache_tag_reg[4][11]  ( .ip(n7173), .ck(clk), .q(\cache_tag[4][11] )
         );
  dp_1 \cache_tag_reg[4][12]  ( .ip(n7155), .ck(clk), .q(\cache_tag[4][12] )
         );
  dp_1 \cache_tag_reg[4][13]  ( .ip(n7137), .ck(clk), .q(\cache_tag[4][13] )
         );
  dp_1 \cache_tag_reg[4][14]  ( .ip(n7119), .ck(clk), .q(\cache_tag[4][14] )
         );
  dp_1 \cache_tag_reg[4][15]  ( .ip(n7101), .ck(clk), .q(\cache_tag[4][15] )
         );
  dp_1 \cache_tag_reg[4][16]  ( .ip(n7083), .ck(clk), .q(\cache_tag[4][16] )
         );
  dp_1 \cache_tag_reg[4][17]  ( .ip(n7065), .ck(clk), .q(\cache_tag[4][17] )
         );
  dp_1 \cache_tag_reg[4][18]  ( .ip(n7047), .ck(clk), .q(\cache_tag[4][18] )
         );
  dp_1 \cache_tag_reg[4][19]  ( .ip(n7029), .ck(clk), .q(\cache_tag[4][19] )
         );
  dp_1 \cache_tag_reg[4][20]  ( .ip(n7011), .ck(clk), .q(\cache_tag[4][20] )
         );
  dp_1 \cache_tag_reg[4][21]  ( .ip(n6993), .ck(clk), .q(\cache_tag[4][21] )
         );
  dp_1 \cache_tag_reg[4][22]  ( .ip(n6975), .ck(clk), .q(\cache_tag[4][22] )
         );
  dp_1 \cache_tag_reg[4][23]  ( .ip(n6957), .ck(clk), .q(\cache_tag[4][23] )
         );
  dp_1 \cache_tag_reg[5][0]  ( .ip(n7370), .ck(clk), .q(\cache_tag[5][0] ) );
  dp_1 \cache_tag_reg[5][1]  ( .ip(n7352), .ck(clk), .q(\cache_tag[5][1] ) );
  dp_1 \cache_tag_reg[5][2]  ( .ip(n7334), .ck(clk), .q(\cache_tag[5][2] ) );
  dp_1 \cache_tag_reg[5][3]  ( .ip(n7316), .ck(clk), .q(\cache_tag[5][3] ) );
  dp_1 \cache_tag_reg[5][4]  ( .ip(n7298), .ck(clk), .q(\cache_tag[5][4] ) );
  dp_1 \cache_tag_reg[5][5]  ( .ip(n7280), .ck(clk), .q(\cache_tag[5][5] ) );
  dp_1 \cache_tag_reg[5][6]  ( .ip(n7262), .ck(clk), .q(\cache_tag[5][6] ) );
  dp_1 \cache_tag_reg[5][7]  ( .ip(n7244), .ck(clk), .q(\cache_tag[5][7] ) );
  dp_1 \cache_tag_reg[5][8]  ( .ip(n7226), .ck(clk), .q(\cache_tag[5][8] ) );
  dp_1 \cache_tag_reg[5][9]  ( .ip(n7208), .ck(clk), .q(\cache_tag[5][9] ) );
  dp_1 \cache_tag_reg[5][10]  ( .ip(n7190), .ck(clk), .q(\cache_tag[5][10] )
         );
  dp_1 \cache_tag_reg[5][11]  ( .ip(n7172), .ck(clk), .q(\cache_tag[5][11] )
         );
  dp_1 \cache_tag_reg[5][12]  ( .ip(n7154), .ck(clk), .q(\cache_tag[5][12] )
         );
  dp_1 \cache_tag_reg[5][13]  ( .ip(n7136), .ck(clk), .q(\cache_tag[5][13] )
         );
  dp_1 \cache_tag_reg[5][14]  ( .ip(n7118), .ck(clk), .q(\cache_tag[5][14] )
         );
  dp_1 \cache_tag_reg[5][15]  ( .ip(n7100), .ck(clk), .q(\cache_tag[5][15] )
         );
  dp_1 \cache_tag_reg[5][16]  ( .ip(n7082), .ck(clk), .q(\cache_tag[5][16] )
         );
  dp_1 \cache_tag_reg[5][17]  ( .ip(n7064), .ck(clk), .q(\cache_tag[5][17] )
         );
  dp_1 \cache_tag_reg[5][18]  ( .ip(n7046), .ck(clk), .q(\cache_tag[5][18] )
         );
  dp_1 \cache_tag_reg[5][19]  ( .ip(n7028), .ck(clk), .q(\cache_tag[5][19] )
         );
  dp_1 \cache_tag_reg[5][20]  ( .ip(n7010), .ck(clk), .q(\cache_tag[5][20] )
         );
  dp_1 \cache_tag_reg[5][21]  ( .ip(n6992), .ck(clk), .q(\cache_tag[5][21] )
         );
  dp_1 \cache_tag_reg[5][22]  ( .ip(n6974), .ck(clk), .q(\cache_tag[5][22] )
         );
  dp_1 \cache_tag_reg[5][23]  ( .ip(n6956), .ck(clk), .q(\cache_tag[5][23] )
         );
  dp_1 \cache_tag_reg[6][0]  ( .ip(n7369), .ck(clk), .q(\cache_tag[6][0] ) );
  dp_1 \cache_tag_reg[6][1]  ( .ip(n7351), .ck(clk), .q(\cache_tag[6][1] ) );
  dp_1 \cache_tag_reg[6][2]  ( .ip(n7333), .ck(clk), .q(\cache_tag[6][2] ) );
  dp_1 \cache_tag_reg[6][3]  ( .ip(n7315), .ck(clk), .q(\cache_tag[6][3] ) );
  dp_1 \cache_tag_reg[6][4]  ( .ip(n7297), .ck(clk), .q(\cache_tag[6][4] ) );
  dp_1 \cache_tag_reg[6][5]  ( .ip(n7279), .ck(clk), .q(\cache_tag[6][5] ) );
  dp_1 \cache_tag_reg[6][6]  ( .ip(n7261), .ck(clk), .q(\cache_tag[6][6] ) );
  dp_1 \cache_tag_reg[6][7]  ( .ip(n7243), .ck(clk), .q(\cache_tag[6][7] ) );
  dp_1 \cache_tag_reg[6][8]  ( .ip(n7225), .ck(clk), .q(\cache_tag[6][8] ) );
  dp_1 \cache_tag_reg[6][9]  ( .ip(n7207), .ck(clk), .q(\cache_tag[6][9] ) );
  dp_1 \cache_tag_reg[6][10]  ( .ip(n7189), .ck(clk), .q(\cache_tag[6][10] )
         );
  dp_1 \cache_tag_reg[6][11]  ( .ip(n7171), .ck(clk), .q(\cache_tag[6][11] )
         );
  dp_1 \cache_tag_reg[6][12]  ( .ip(n7153), .ck(clk), .q(\cache_tag[6][12] )
         );
  dp_1 \cache_tag_reg[6][13]  ( .ip(n7135), .ck(clk), .q(\cache_tag[6][13] )
         );
  dp_1 \cache_tag_reg[6][14]  ( .ip(n7117), .ck(clk), .q(\cache_tag[6][14] )
         );
  dp_1 \cache_tag_reg[6][15]  ( .ip(n7099), .ck(clk), .q(\cache_tag[6][15] )
         );
  dp_1 \cache_tag_reg[6][16]  ( .ip(n7081), .ck(clk), .q(\cache_tag[6][16] )
         );
  dp_1 \cache_tag_reg[6][17]  ( .ip(n7063), .ck(clk), .q(\cache_tag[6][17] )
         );
  dp_1 \cache_tag_reg[6][18]  ( .ip(n7045), .ck(clk), .q(\cache_tag[6][18] )
         );
  dp_1 \cache_tag_reg[6][19]  ( .ip(n7027), .ck(clk), .q(\cache_tag[6][19] )
         );
  dp_1 \cache_tag_reg[6][20]  ( .ip(n7009), .ck(clk), .q(\cache_tag[6][20] )
         );
  dp_1 \cache_tag_reg[6][21]  ( .ip(n6991), .ck(clk), .q(\cache_tag[6][21] )
         );
  dp_1 \cache_tag_reg[6][22]  ( .ip(n6973), .ck(clk), .q(\cache_tag[6][22] )
         );
  dp_1 \cache_tag_reg[6][23]  ( .ip(n6955), .ck(clk), .q(\cache_tag[6][23] )
         );
  dp_1 \cache_tag_reg[7][0]  ( .ip(n7368), .ck(clk), .q(\cache_tag[7][0] ) );
  dp_1 \cache_tag_reg[7][1]  ( .ip(n7350), .ck(clk), .q(\cache_tag[7][1] ) );
  dp_1 \cache_tag_reg[7][2]  ( .ip(n7332), .ck(clk), .q(\cache_tag[7][2] ) );
  dp_1 \cache_tag_reg[7][3]  ( .ip(n7314), .ck(clk), .q(\cache_tag[7][3] ) );
  dp_1 \cache_tag_reg[7][4]  ( .ip(n7296), .ck(clk), .q(\cache_tag[7][4] ) );
  dp_1 \cache_tag_reg[7][5]  ( .ip(n7278), .ck(clk), .q(\cache_tag[7][5] ) );
  dp_1 \cache_tag_reg[7][6]  ( .ip(n7260), .ck(clk), .q(\cache_tag[7][6] ) );
  dp_1 \cache_tag_reg[7][7]  ( .ip(n7242), .ck(clk), .q(\cache_tag[7][7] ) );
  dp_1 \cache_tag_reg[7][8]  ( .ip(n7224), .ck(clk), .q(\cache_tag[7][8] ) );
  dp_1 \cache_tag_reg[7][9]  ( .ip(n7206), .ck(clk), .q(\cache_tag[7][9] ) );
  dp_1 \cache_tag_reg[7][10]  ( .ip(n7188), .ck(clk), .q(\cache_tag[7][10] )
         );
  dp_1 \cache_tag_reg[7][11]  ( .ip(n7170), .ck(clk), .q(\cache_tag[7][11] )
         );
  dp_1 \cache_tag_reg[7][12]  ( .ip(n7152), .ck(clk), .q(\cache_tag[7][12] )
         );
  dp_1 \cache_tag_reg[7][13]  ( .ip(n7134), .ck(clk), .q(\cache_tag[7][13] )
         );
  dp_1 \cache_tag_reg[7][14]  ( .ip(n7116), .ck(clk), .q(\cache_tag[7][14] )
         );
  dp_1 \cache_tag_reg[7][15]  ( .ip(n7098), .ck(clk), .q(\cache_tag[7][15] )
         );
  dp_1 \cache_tag_reg[7][16]  ( .ip(n7080), .ck(clk), .q(\cache_tag[7][16] )
         );
  dp_1 \cache_tag_reg[7][17]  ( .ip(n7062), .ck(clk), .q(\cache_tag[7][17] )
         );
  dp_1 \cache_tag_reg[7][18]  ( .ip(n7044), .ck(clk), .q(\cache_tag[7][18] )
         );
  dp_1 \cache_tag_reg[7][19]  ( .ip(n7026), .ck(clk), .q(\cache_tag[7][19] )
         );
  dp_1 \cache_tag_reg[7][20]  ( .ip(n7008), .ck(clk), .q(\cache_tag[7][20] )
         );
  dp_1 \cache_tag_reg[7][21]  ( .ip(n6990), .ck(clk), .q(\cache_tag[7][21] )
         );
  dp_1 \cache_tag_reg[7][22]  ( .ip(n6972), .ck(clk), .q(\cache_tag[7][22] )
         );
  dp_1 \cache_tag_reg[7][23]  ( .ip(n6954), .ck(clk), .q(\cache_tag[7][23] )
         );
  dp_1 \cache_tag_reg[8][0]  ( .ip(n7367), .ck(clk), .q(\cache_tag[8][0] ) );
  dp_1 \cache_tag_reg[8][1]  ( .ip(n7349), .ck(clk), .q(\cache_tag[8][1] ) );
  dp_1 \cache_tag_reg[8][2]  ( .ip(n7331), .ck(clk), .q(\cache_tag[8][2] ) );
  dp_1 \cache_tag_reg[8][3]  ( .ip(n7313), .ck(clk), .q(\cache_tag[8][3] ) );
  dp_1 \cache_tag_reg[8][4]  ( .ip(n7295), .ck(clk), .q(\cache_tag[8][4] ) );
  dp_1 \cache_tag_reg[8][5]  ( .ip(n7277), .ck(clk), .q(\cache_tag[8][5] ) );
  dp_1 \cache_tag_reg[8][6]  ( .ip(n7259), .ck(clk), .q(\cache_tag[8][6] ) );
  dp_1 \cache_tag_reg[8][7]  ( .ip(n7241), .ck(clk), .q(\cache_tag[8][7] ) );
  dp_1 \cache_tag_reg[8][8]  ( .ip(n7223), .ck(clk), .q(\cache_tag[8][8] ) );
  dp_1 \cache_tag_reg[8][9]  ( .ip(n7205), .ck(clk), .q(\cache_tag[8][9] ) );
  dp_1 \cache_tag_reg[8][10]  ( .ip(n7187), .ck(clk), .q(\cache_tag[8][10] )
         );
  dp_1 \cache_tag_reg[8][11]  ( .ip(n7169), .ck(clk), .q(\cache_tag[8][11] )
         );
  dp_1 \cache_tag_reg[8][12]  ( .ip(n7151), .ck(clk), .q(\cache_tag[8][12] )
         );
  dp_1 \cache_tag_reg[8][13]  ( .ip(n7133), .ck(clk), .q(\cache_tag[8][13] )
         );
  dp_1 \cache_tag_reg[8][14]  ( .ip(n7115), .ck(clk), .q(\cache_tag[8][14] )
         );
  dp_1 \cache_tag_reg[8][15]  ( .ip(n7097), .ck(clk), .q(\cache_tag[8][15] )
         );
  dp_1 \cache_tag_reg[8][16]  ( .ip(n7079), .ck(clk), .q(\cache_tag[8][16] )
         );
  dp_1 \cache_tag_reg[8][17]  ( .ip(n7061), .ck(clk), .q(\cache_tag[8][17] )
         );
  dp_1 \cache_tag_reg[8][18]  ( .ip(n7043), .ck(clk), .q(\cache_tag[8][18] )
         );
  dp_1 \cache_tag_reg[8][19]  ( .ip(n7025), .ck(clk), .q(\cache_tag[8][19] )
         );
  dp_1 \cache_tag_reg[8][20]  ( .ip(n7007), .ck(clk), .q(\cache_tag[8][20] )
         );
  dp_1 \cache_tag_reg[8][21]  ( .ip(n6989), .ck(clk), .q(\cache_tag[8][21] )
         );
  dp_1 \cache_tag_reg[8][22]  ( .ip(n6971), .ck(clk), .q(\cache_tag[8][22] )
         );
  dp_1 \cache_tag_reg[8][23]  ( .ip(n6953), .ck(clk), .q(\cache_tag[8][23] )
         );
  dp_1 \cache_tag_reg[9][0]  ( .ip(n7366), .ck(clk), .q(\cache_tag[9][0] ) );
  dp_1 \cache_tag_reg[9][1]  ( .ip(n7348), .ck(clk), .q(\cache_tag[9][1] ) );
  dp_1 \cache_tag_reg[9][2]  ( .ip(n7330), .ck(clk), .q(\cache_tag[9][2] ) );
  dp_1 \cache_tag_reg[9][3]  ( .ip(n7312), .ck(clk), .q(\cache_tag[9][3] ) );
  dp_1 \cache_tag_reg[9][4]  ( .ip(n7294), .ck(clk), .q(\cache_tag[9][4] ) );
  dp_1 \cache_tag_reg[9][5]  ( .ip(n7276), .ck(clk), .q(\cache_tag[9][5] ) );
  dp_1 \cache_tag_reg[9][6]  ( .ip(n7258), .ck(clk), .q(\cache_tag[9][6] ) );
  dp_1 \cache_tag_reg[9][7]  ( .ip(n7240), .ck(clk), .q(\cache_tag[9][7] ) );
  dp_1 \cache_tag_reg[9][8]  ( .ip(n7222), .ck(clk), .q(\cache_tag[9][8] ) );
  dp_1 \cache_tag_reg[9][9]  ( .ip(n7204), .ck(clk), .q(\cache_tag[9][9] ) );
  dp_1 \cache_tag_reg[9][10]  ( .ip(n7186), .ck(clk), .q(\cache_tag[9][10] )
         );
  dp_1 \cache_tag_reg[9][11]  ( .ip(n7168), .ck(clk), .q(\cache_tag[9][11] )
         );
  dp_1 \cache_tag_reg[9][12]  ( .ip(n7150), .ck(clk), .q(\cache_tag[9][12] )
         );
  dp_1 \cache_tag_reg[9][13]  ( .ip(n7132), .ck(clk), .q(\cache_tag[9][13] )
         );
  dp_1 \cache_tag_reg[9][14]  ( .ip(n7114), .ck(clk), .q(\cache_tag[9][14] )
         );
  dp_1 \cache_tag_reg[9][15]  ( .ip(n7096), .ck(clk), .q(\cache_tag[9][15] )
         );
  dp_1 \cache_tag_reg[9][16]  ( .ip(n7078), .ck(clk), .q(\cache_tag[9][16] )
         );
  dp_1 \cache_tag_reg[9][17]  ( .ip(n7060), .ck(clk), .q(\cache_tag[9][17] )
         );
  dp_1 \cache_tag_reg[9][18]  ( .ip(n7042), .ck(clk), .q(\cache_tag[9][18] )
         );
  dp_1 \cache_tag_reg[9][19]  ( .ip(n7024), .ck(clk), .q(\cache_tag[9][19] )
         );
  dp_1 \cache_tag_reg[9][20]  ( .ip(n7006), .ck(clk), .q(\cache_tag[9][20] )
         );
  dp_1 \cache_tag_reg[9][21]  ( .ip(n6988), .ck(clk), .q(\cache_tag[9][21] )
         );
  dp_1 \cache_tag_reg[9][22]  ( .ip(n6970), .ck(clk), .q(\cache_tag[9][22] )
         );
  dp_1 \cache_tag_reg[9][23]  ( .ip(n6952), .ck(clk), .q(\cache_tag[9][23] )
         );
  dp_1 \cache_tag_reg[10][0]  ( .ip(n7365), .ck(clk), .q(\cache_tag[10][0] )
         );
  dp_1 \cache_tag_reg[10][1]  ( .ip(n7347), .ck(clk), .q(\cache_tag[10][1] )
         );
  dp_1 \cache_tag_reg[10][2]  ( .ip(n7329), .ck(clk), .q(\cache_tag[10][2] )
         );
  dp_1 \cache_tag_reg[10][3]  ( .ip(n7311), .ck(clk), .q(\cache_tag[10][3] )
         );
  dp_1 \cache_tag_reg[10][4]  ( .ip(n7293), .ck(clk), .q(\cache_tag[10][4] )
         );
  dp_1 \cache_tag_reg[10][5]  ( .ip(n7275), .ck(clk), .q(\cache_tag[10][5] )
         );
  dp_1 \cache_tag_reg[10][6]  ( .ip(n7257), .ck(clk), .q(\cache_tag[10][6] )
         );
  dp_1 \cache_tag_reg[10][7]  ( .ip(n7239), .ck(clk), .q(\cache_tag[10][7] )
         );
  dp_1 \cache_tag_reg[10][8]  ( .ip(n7221), .ck(clk), .q(\cache_tag[10][8] )
         );
  dp_1 \cache_tag_reg[10][9]  ( .ip(n7203), .ck(clk), .q(\cache_tag[10][9] )
         );
  dp_1 \cache_tag_reg[10][10]  ( .ip(n7185), .ck(clk), .q(\cache_tag[10][10] )
         );
  dp_1 \cache_tag_reg[10][11]  ( .ip(n7167), .ck(clk), .q(\cache_tag[10][11] )
         );
  dp_1 \cache_tag_reg[10][12]  ( .ip(n7149), .ck(clk), .q(\cache_tag[10][12] )
         );
  dp_1 \cache_tag_reg[10][13]  ( .ip(n7131), .ck(clk), .q(\cache_tag[10][13] )
         );
  dp_1 \cache_tag_reg[10][14]  ( .ip(n7113), .ck(clk), .q(\cache_tag[10][14] )
         );
  dp_1 \cache_tag_reg[10][15]  ( .ip(n7095), .ck(clk), .q(\cache_tag[10][15] )
         );
  dp_1 \cache_tag_reg[10][16]  ( .ip(n7077), .ck(clk), .q(\cache_tag[10][16] )
         );
  dp_1 \cache_tag_reg[10][17]  ( .ip(n7059), .ck(clk), .q(\cache_tag[10][17] )
         );
  dp_1 \cache_tag_reg[10][18]  ( .ip(n7041), .ck(clk), .q(\cache_tag[10][18] )
         );
  dp_1 \cache_tag_reg[10][19]  ( .ip(n7023), .ck(clk), .q(\cache_tag[10][19] )
         );
  dp_1 \cache_tag_reg[10][20]  ( .ip(n7005), .ck(clk), .q(\cache_tag[10][20] )
         );
  dp_1 \cache_tag_reg[10][21]  ( .ip(n6987), .ck(clk), .q(\cache_tag[10][21] )
         );
  dp_1 \cache_tag_reg[10][22]  ( .ip(n6969), .ck(clk), .q(\cache_tag[10][22] )
         );
  dp_1 \cache_tag_reg[10][23]  ( .ip(n6951), .ck(clk), .q(\cache_tag[10][23] )
         );
  dp_1 \cache_tag_reg[11][0]  ( .ip(n7364), .ck(clk), .q(\cache_tag[11][0] )
         );
  dp_1 \cache_tag_reg[11][1]  ( .ip(n7346), .ck(clk), .q(\cache_tag[11][1] )
         );
  dp_1 \cache_tag_reg[11][2]  ( .ip(n7328), .ck(clk), .q(\cache_tag[11][2] )
         );
  dp_1 \cache_tag_reg[11][3]  ( .ip(n7310), .ck(clk), .q(\cache_tag[11][3] )
         );
  dp_1 \cache_tag_reg[11][4]  ( .ip(n7292), .ck(clk), .q(\cache_tag[11][4] )
         );
  dp_1 \cache_tag_reg[11][5]  ( .ip(n7274), .ck(clk), .q(\cache_tag[11][5] )
         );
  dp_1 \cache_tag_reg[11][6]  ( .ip(n7256), .ck(clk), .q(\cache_tag[11][6] )
         );
  dp_1 \cache_tag_reg[11][7]  ( .ip(n7238), .ck(clk), .q(\cache_tag[11][7] )
         );
  dp_1 \cache_tag_reg[11][8]  ( .ip(n7220), .ck(clk), .q(\cache_tag[11][8] )
         );
  dp_1 \cache_tag_reg[11][9]  ( .ip(n7202), .ck(clk), .q(\cache_tag[11][9] )
         );
  dp_1 \cache_tag_reg[11][10]  ( .ip(n7184), .ck(clk), .q(\cache_tag[11][10] )
         );
  dp_1 \cache_tag_reg[11][11]  ( .ip(n7166), .ck(clk), .q(\cache_tag[11][11] )
         );
  dp_1 \cache_tag_reg[11][12]  ( .ip(n7148), .ck(clk), .q(\cache_tag[11][12] )
         );
  dp_1 \cache_tag_reg[11][13]  ( .ip(n7130), .ck(clk), .q(\cache_tag[11][13] )
         );
  dp_1 \cache_tag_reg[11][14]  ( .ip(n7112), .ck(clk), .q(\cache_tag[11][14] )
         );
  dp_1 \cache_tag_reg[11][15]  ( .ip(n7094), .ck(clk), .q(\cache_tag[11][15] )
         );
  dp_1 \cache_tag_reg[11][16]  ( .ip(n7076), .ck(clk), .q(\cache_tag[11][16] )
         );
  dp_1 \cache_tag_reg[11][17]  ( .ip(n7058), .ck(clk), .q(\cache_tag[11][17] )
         );
  dp_1 \cache_tag_reg[11][18]  ( .ip(n7040), .ck(clk), .q(\cache_tag[11][18] )
         );
  dp_1 \cache_tag_reg[11][19]  ( .ip(n7022), .ck(clk), .q(\cache_tag[11][19] )
         );
  dp_1 \cache_tag_reg[11][20]  ( .ip(n7004), .ck(clk), .q(\cache_tag[11][20] )
         );
  dp_1 \cache_tag_reg[11][21]  ( .ip(n6986), .ck(clk), .q(\cache_tag[11][21] )
         );
  dp_1 \cache_tag_reg[11][22]  ( .ip(n6968), .ck(clk), .q(\cache_tag[11][22] )
         );
  dp_1 \cache_tag_reg[11][23]  ( .ip(n6950), .ck(clk), .q(\cache_tag[11][23] )
         );
  dp_1 \cache_tag_reg[12][0]  ( .ip(n7363), .ck(clk), .q(\cache_tag[12][0] )
         );
  dp_1 \cache_tag_reg[12][1]  ( .ip(n7345), .ck(clk), .q(\cache_tag[12][1] )
         );
  dp_1 \cache_tag_reg[12][2]  ( .ip(n7327), .ck(clk), .q(\cache_tag[12][2] )
         );
  dp_1 \cache_tag_reg[12][3]  ( .ip(n7309), .ck(clk), .q(\cache_tag[12][3] )
         );
  dp_1 \cache_tag_reg[12][4]  ( .ip(n7291), .ck(clk), .q(\cache_tag[12][4] )
         );
  dp_1 \cache_tag_reg[12][5]  ( .ip(n7273), .ck(clk), .q(\cache_tag[12][5] )
         );
  dp_1 \cache_tag_reg[12][6]  ( .ip(n7255), .ck(clk), .q(\cache_tag[12][6] )
         );
  dp_1 \cache_tag_reg[12][7]  ( .ip(n7237), .ck(clk), .q(\cache_tag[12][7] )
         );
  dp_1 \cache_tag_reg[12][8]  ( .ip(n7219), .ck(clk), .q(\cache_tag[12][8] )
         );
  dp_1 \cache_tag_reg[12][9]  ( .ip(n7201), .ck(clk), .q(\cache_tag[12][9] )
         );
  dp_1 \cache_tag_reg[12][10]  ( .ip(n7183), .ck(clk), .q(\cache_tag[12][10] )
         );
  dp_1 \cache_tag_reg[12][11]  ( .ip(n7165), .ck(clk), .q(\cache_tag[12][11] )
         );
  dp_1 \cache_tag_reg[12][12]  ( .ip(n7147), .ck(clk), .q(\cache_tag[12][12] )
         );
  dp_1 \cache_tag_reg[12][13]  ( .ip(n7129), .ck(clk), .q(\cache_tag[12][13] )
         );
  dp_1 \cache_tag_reg[12][14]  ( .ip(n7111), .ck(clk), .q(\cache_tag[12][14] )
         );
  dp_1 \cache_tag_reg[12][15]  ( .ip(n7093), .ck(clk), .q(\cache_tag[12][15] )
         );
  dp_1 \cache_tag_reg[12][16]  ( .ip(n7075), .ck(clk), .q(\cache_tag[12][16] )
         );
  dp_1 \cache_tag_reg[12][17]  ( .ip(n7057), .ck(clk), .q(\cache_tag[12][17] )
         );
  dp_1 \cache_tag_reg[12][18]  ( .ip(n7039), .ck(clk), .q(\cache_tag[12][18] )
         );
  dp_1 \cache_tag_reg[12][19]  ( .ip(n7021), .ck(clk), .q(\cache_tag[12][19] )
         );
  dp_1 \cache_tag_reg[12][20]  ( .ip(n7003), .ck(clk), .q(\cache_tag[12][20] )
         );
  dp_1 \cache_tag_reg[12][21]  ( .ip(n6985), .ck(clk), .q(\cache_tag[12][21] )
         );
  dp_1 \cache_tag_reg[12][22]  ( .ip(n6967), .ck(clk), .q(\cache_tag[12][22] )
         );
  dp_1 \cache_tag_reg[12][23]  ( .ip(n6949), .ck(clk), .q(\cache_tag[12][23] )
         );
  dp_1 \cache_tag_reg[13][0]  ( .ip(n7362), .ck(clk), .q(\cache_tag[13][0] )
         );
  dp_1 \cache_tag_reg[13][1]  ( .ip(n7344), .ck(clk), .q(\cache_tag[13][1] )
         );
  dp_1 \cache_tag_reg[13][2]  ( .ip(n7326), .ck(clk), .q(\cache_tag[13][2] )
         );
  dp_1 \cache_tag_reg[13][3]  ( .ip(n7308), .ck(clk), .q(\cache_tag[13][3] )
         );
  dp_1 \cache_tag_reg[13][4]  ( .ip(n7290), .ck(clk), .q(\cache_tag[13][4] )
         );
  dp_1 \cache_tag_reg[13][5]  ( .ip(n7272), .ck(clk), .q(\cache_tag[13][5] )
         );
  dp_1 \cache_tag_reg[13][6]  ( .ip(n7254), .ck(clk), .q(\cache_tag[13][6] )
         );
  dp_1 \cache_tag_reg[13][7]  ( .ip(n7236), .ck(clk), .q(\cache_tag[13][7] )
         );
  dp_1 \cache_tag_reg[13][8]  ( .ip(n7218), .ck(clk), .q(\cache_tag[13][8] )
         );
  dp_1 \cache_tag_reg[13][9]  ( .ip(n7200), .ck(clk), .q(\cache_tag[13][9] )
         );
  dp_1 \cache_tag_reg[13][10]  ( .ip(n7182), .ck(clk), .q(\cache_tag[13][10] )
         );
  dp_1 \cache_tag_reg[13][11]  ( .ip(n7164), .ck(clk), .q(\cache_tag[13][11] )
         );
  dp_1 \cache_tag_reg[13][12]  ( .ip(n7146), .ck(clk), .q(\cache_tag[13][12] )
         );
  dp_1 \cache_tag_reg[13][13]  ( .ip(n7128), .ck(clk), .q(\cache_tag[13][13] )
         );
  dp_1 \cache_tag_reg[13][14]  ( .ip(n7110), .ck(clk), .q(\cache_tag[13][14] )
         );
  dp_1 \cache_tag_reg[13][15]  ( .ip(n7092), .ck(clk), .q(\cache_tag[13][15] )
         );
  dp_1 \cache_tag_reg[13][16]  ( .ip(n7074), .ck(clk), .q(\cache_tag[13][16] )
         );
  dp_1 \cache_tag_reg[13][17]  ( .ip(n7056), .ck(clk), .q(\cache_tag[13][17] )
         );
  dp_1 \cache_tag_reg[13][18]  ( .ip(n7038), .ck(clk), .q(\cache_tag[13][18] )
         );
  dp_1 \cache_tag_reg[13][19]  ( .ip(n7020), .ck(clk), .q(\cache_tag[13][19] )
         );
  dp_1 \cache_tag_reg[13][20]  ( .ip(n7002), .ck(clk), .q(\cache_tag[13][20] )
         );
  dp_1 \cache_tag_reg[13][21]  ( .ip(n6984), .ck(clk), .q(\cache_tag[13][21] )
         );
  dp_1 \cache_tag_reg[13][22]  ( .ip(n6966), .ck(clk), .q(\cache_tag[13][22] )
         );
  dp_1 \cache_tag_reg[13][23]  ( .ip(n6948), .ck(clk), .q(\cache_tag[13][23] )
         );
  dp_1 \cache_tag_reg[14][0]  ( .ip(n7361), .ck(clk), .q(\cache_tag[14][0] )
         );
  dp_1 \cache_tag_reg[14][1]  ( .ip(n7343), .ck(clk), .q(\cache_tag[14][1] )
         );
  dp_1 \cache_tag_reg[14][2]  ( .ip(n7325), .ck(clk), .q(\cache_tag[14][2] )
         );
  dp_1 \cache_tag_reg[14][3]  ( .ip(n7307), .ck(clk), .q(\cache_tag[14][3] )
         );
  dp_1 \cache_tag_reg[14][4]  ( .ip(n7289), .ck(clk), .q(\cache_tag[14][4] )
         );
  dp_1 \cache_tag_reg[14][5]  ( .ip(n7271), .ck(clk), .q(\cache_tag[14][5] )
         );
  dp_1 \cache_tag_reg[14][6]  ( .ip(n7253), .ck(clk), .q(\cache_tag[14][6] )
         );
  dp_1 \cache_tag_reg[14][7]  ( .ip(n7235), .ck(clk), .q(\cache_tag[14][7] )
         );
  dp_1 \cache_tag_reg[14][8]  ( .ip(n7217), .ck(clk), .q(\cache_tag[14][8] )
         );
  dp_1 \cache_tag_reg[14][9]  ( .ip(n7199), .ck(clk), .q(\cache_tag[14][9] )
         );
  dp_1 \cache_tag_reg[14][10]  ( .ip(n7181), .ck(clk), .q(\cache_tag[14][10] )
         );
  dp_1 \cache_tag_reg[14][11]  ( .ip(n7163), .ck(clk), .q(\cache_tag[14][11] )
         );
  dp_1 \cache_tag_reg[14][12]  ( .ip(n7145), .ck(clk), .q(\cache_tag[14][12] )
         );
  dp_1 \cache_tag_reg[14][13]  ( .ip(n7127), .ck(clk), .q(\cache_tag[14][13] )
         );
  dp_1 \cache_tag_reg[14][14]  ( .ip(n7109), .ck(clk), .q(\cache_tag[14][14] )
         );
  dp_1 \cache_tag_reg[14][15]  ( .ip(n7091), .ck(clk), .q(\cache_tag[14][15] )
         );
  dp_1 \cache_tag_reg[14][16]  ( .ip(n7073), .ck(clk), .q(\cache_tag[14][16] )
         );
  dp_1 \cache_tag_reg[14][17]  ( .ip(n7055), .ck(clk), .q(\cache_tag[14][17] )
         );
  dp_1 \cache_tag_reg[14][18]  ( .ip(n7037), .ck(clk), .q(\cache_tag[14][18] )
         );
  dp_1 \cache_tag_reg[14][19]  ( .ip(n7019), .ck(clk), .q(\cache_tag[14][19] )
         );
  dp_1 \cache_tag_reg[14][20]  ( .ip(n7001), .ck(clk), .q(\cache_tag[14][20] )
         );
  dp_1 \cache_tag_reg[14][21]  ( .ip(n6983), .ck(clk), .q(\cache_tag[14][21] )
         );
  dp_1 \cache_tag_reg[14][22]  ( .ip(n6965), .ck(clk), .q(\cache_tag[14][22] )
         );
  dp_1 \cache_tag_reg[14][23]  ( .ip(n6947), .ck(clk), .q(\cache_tag[14][23] )
         );
  dp_1 \cache_tag_reg[15][0]  ( .ip(n7360), .ck(clk), .q(\cache_tag[15][0] )
         );
  dp_1 \cache_tag_reg[15][1]  ( .ip(n7342), .ck(clk), .q(\cache_tag[15][1] )
         );
  dp_1 \cache_tag_reg[15][2]  ( .ip(n7324), .ck(clk), .q(\cache_tag[15][2] )
         );
  dp_1 \cache_tag_reg[15][3]  ( .ip(n7306), .ck(clk), .q(\cache_tag[15][3] )
         );
  dp_1 \cache_tag_reg[15][4]  ( .ip(n7288), .ck(clk), .q(\cache_tag[15][4] )
         );
  dp_1 \cache_tag_reg[15][5]  ( .ip(n7270), .ck(clk), .q(\cache_tag[15][5] )
         );
  dp_1 \cache_tag_reg[15][6]  ( .ip(n7252), .ck(clk), .q(\cache_tag[15][6] )
         );
  dp_1 \cache_tag_reg[15][7]  ( .ip(n7234), .ck(clk), .q(\cache_tag[15][7] )
         );
  dp_1 \cache_tag_reg[15][8]  ( .ip(n7216), .ck(clk), .q(\cache_tag[15][8] )
         );
  dp_1 \cache_tag_reg[15][9]  ( .ip(n7198), .ck(clk), .q(\cache_tag[15][9] )
         );
  dp_1 \cache_tag_reg[15][10]  ( .ip(n7180), .ck(clk), .q(\cache_tag[15][10] )
         );
  dp_1 \cache_tag_reg[15][11]  ( .ip(n7162), .ck(clk), .q(\cache_tag[15][11] )
         );
  dp_1 \cache_tag_reg[15][12]  ( .ip(n7144), .ck(clk), .q(\cache_tag[15][12] )
         );
  dp_1 \cache_tag_reg[15][13]  ( .ip(n7126), .ck(clk), .q(\cache_tag[15][13] )
         );
  dp_1 \cache_tag_reg[15][14]  ( .ip(n7108), .ck(clk), .q(\cache_tag[15][14] )
         );
  dp_1 \cache_tag_reg[15][15]  ( .ip(n7090), .ck(clk), .q(\cache_tag[15][15] )
         );
  dp_1 \cache_tag_reg[15][16]  ( .ip(n7072), .ck(clk), .q(\cache_tag[15][16] )
         );
  dp_1 \cache_tag_reg[15][17]  ( .ip(n7054), .ck(clk), .q(\cache_tag[15][17] )
         );
  dp_1 \cache_tag_reg[15][18]  ( .ip(n7036), .ck(clk), .q(\cache_tag[15][18] )
         );
  dp_1 \cache_tag_reg[15][19]  ( .ip(n7018), .ck(clk), .q(\cache_tag[15][19] )
         );
  dp_1 \cache_tag_reg[15][20]  ( .ip(n7000), .ck(clk), .q(\cache_tag[15][20] )
         );
  dp_1 \cache_tag_reg[15][21]  ( .ip(n6982), .ck(clk), .q(\cache_tag[15][21] )
         );
  dp_1 \cache_tag_reg[15][22]  ( .ip(n6964), .ck(clk), .q(\cache_tag[15][22] )
         );
  dp_1 \cache_tag_reg[15][23]  ( .ip(n6946), .ck(clk), .q(\cache_tag[15][23] )
         );
  dp_1 \data_rd_reg[0]  ( .ip(n6944), .ck(clk), .q(N3519) );
  dp_1 \data_rd_reg[1]  ( .ip(n6942), .ck(clk), .q(N3516) );
  dp_1 \data_rd_reg[2]  ( .ip(n6940), .ck(clk), .q(N3513) );
  dp_1 \data_rd_reg[3]  ( .ip(n6938), .ck(clk), .q(N3510) );
  dp_1 \data_rd_reg[4]  ( .ip(n6936), .ck(clk), .q(N3507) );
  dp_1 \data_rd_reg[5]  ( .ip(n6934), .ck(clk), .q(N3504) );
  dp_1 \data_rd_reg[6]  ( .ip(n6932), .ck(clk), .q(N3501) );
  dp_1 \data_rd_reg[7]  ( .ip(n6930), .ck(clk), .q(N3498) );
  dp_1 \data_rd_reg[8]  ( .ip(n6928), .ck(clk), .q(N3495) );
  dp_1 \data_rd_reg[9]  ( .ip(n6926), .ck(clk), .q(N3492) );
  dp_1 \data_rd_reg[10]  ( .ip(n6924), .ck(clk), .q(N3489) );
  dp_1 \data_rd_reg[11]  ( .ip(n6922), .ck(clk), .q(N3486) );
  dp_1 \data_rd_reg[12]  ( .ip(n6920), .ck(clk), .q(N3483) );
  dp_1 \data_rd_reg[13]  ( .ip(n6918), .ck(clk), .q(N3480) );
  dp_1 \data_rd_reg[14]  ( .ip(n6916), .ck(clk), .q(N3477) );
  dp_1 \data_rd_reg[15]  ( .ip(n6914), .ck(clk), .q(N3474) );
  dp_1 \data_rd_reg[16]  ( .ip(n6912), .ck(clk), .q(N3471) );
  dp_1 \data_rd_reg[17]  ( .ip(n6910), .ck(clk), .q(N3468) );
  dp_1 \data_rd_reg[18]  ( .ip(n6908), .ck(clk), .q(N3465) );
  dp_1 \data_rd_reg[19]  ( .ip(n6906), .ck(clk), .q(N3462) );
  dp_1 \data_rd_reg[20]  ( .ip(n6904), .ck(clk), .q(N3459) );
  dp_1 \data_rd_reg[21]  ( .ip(n6902), .ck(clk), .q(N3456) );
  dp_1 \data_rd_reg[22]  ( .ip(n6900), .ck(clk), .q(N3453) );
  dp_1 \data_rd_reg[23]  ( .ip(n6898), .ck(clk), .q(N3450) );
  dp_1 \data_rd_reg[24]  ( .ip(n6896), .ck(clk), .q(N3447) );
  dp_1 \data_rd_reg[25]  ( .ip(n6894), .ck(clk), .q(N3444) );
  dp_1 \data_rd_reg[26]  ( .ip(n6892), .ck(clk), .q(N3441) );
  dp_1 \data_rd_reg[27]  ( .ip(n6890), .ck(clk), .q(N3438) );
  dp_1 \data_rd_reg[28]  ( .ip(n6888), .ck(clk), .q(N3435) );
  dp_1 \data_rd_reg[29]  ( .ip(n6886), .ck(clk), .q(N3432) );
  dp_1 \data_rd_reg[30]  ( .ip(n6884), .ck(clk), .q(N3429) );
  dp_1 \data_rd_reg[31]  ( .ip(n6882), .ck(clk), .q(N3426) );
  dp_1 \iCache_data_wr_reg[0]  ( .ip(n6863), .ck(clk), .q(iCache_data_wr[0])
         );
  dp_1 \cache_data_reg[0][0]  ( .ip(n6831), .ck(clk), .q(\cache_data[0][0] )
         );
  dp_1 \cache_data_reg[0][32]  ( .ip(n6799), .ck(clk), .q(\cache_data[0][32] )
         );
  dp_1 \cache_data_reg[0][64]  ( .ip(n6767), .ck(clk), .q(\cache_data[0][64] )
         );
  dp_1 \cache_data_reg[0][96]  ( .ip(n6735), .ck(clk), .q(\cache_data[0][96] )
         );
  dp_1 \cache_data_reg[1][0]  ( .ip(n6703), .ck(clk), .q(\cache_data[1][0] )
         );
  dp_1 \cache_data_reg[1][32]  ( .ip(n6671), .ck(clk), .q(\cache_data[1][32] )
         );
  dp_1 \cache_data_reg[1][64]  ( .ip(n6639), .ck(clk), .q(\cache_data[1][64] )
         );
  dp_1 \cache_data_reg[1][96]  ( .ip(n6607), .ck(clk), .q(\cache_data[1][96] )
         );
  dp_1 \cache_data_reg[2][0]  ( .ip(n6575), .ck(clk), .q(\cache_data[2][0] )
         );
  dp_1 \cache_data_reg[2][32]  ( .ip(n6543), .ck(clk), .q(\cache_data[2][32] )
         );
  dp_1 \cache_data_reg[2][64]  ( .ip(n6511), .ck(clk), .q(\cache_data[2][64] )
         );
  dp_1 \cache_data_reg[2][96]  ( .ip(n6479), .ck(clk), .q(\cache_data[2][96] )
         );
  dp_1 \cache_data_reg[3][0]  ( .ip(n6447), .ck(clk), .q(\cache_data[3][0] )
         );
  dp_1 \cache_data_reg[3][32]  ( .ip(n6415), .ck(clk), .q(\cache_data[3][32] )
         );
  dp_1 \cache_data_reg[3][64]  ( .ip(n6383), .ck(clk), .q(\cache_data[3][64] )
         );
  dp_1 \cache_data_reg[3][96]  ( .ip(n6351), .ck(clk), .q(\cache_data[3][96] )
         );
  dp_1 \cache_data_reg[4][0]  ( .ip(n6319), .ck(clk), .q(\cache_data[4][0] )
         );
  dp_1 \cache_data_reg[4][32]  ( .ip(n6287), .ck(clk), .q(\cache_data[4][32] )
         );
  dp_1 \cache_data_reg[4][64]  ( .ip(n6255), .ck(clk), .q(\cache_data[4][64] )
         );
  dp_1 \cache_data_reg[4][96]  ( .ip(n6223), .ck(clk), .q(\cache_data[4][96] )
         );
  dp_1 \cache_data_reg[5][0]  ( .ip(n6191), .ck(clk), .q(\cache_data[5][0] )
         );
  dp_1 \cache_data_reg[5][32]  ( .ip(n6159), .ck(clk), .q(\cache_data[5][32] )
         );
  dp_1 \cache_data_reg[5][64]  ( .ip(n6127), .ck(clk), .q(\cache_data[5][64] )
         );
  dp_1 \cache_data_reg[5][96]  ( .ip(n6095), .ck(clk), .q(\cache_data[5][96] )
         );
  dp_1 \cache_data_reg[6][0]  ( .ip(n6063), .ck(clk), .q(\cache_data[6][0] )
         );
  dp_1 \cache_data_reg[6][32]  ( .ip(n6031), .ck(clk), .q(\cache_data[6][32] )
         );
  dp_1 \cache_data_reg[6][64]  ( .ip(n5999), .ck(clk), .q(\cache_data[6][64] )
         );
  dp_1 \cache_data_reg[6][96]  ( .ip(n5967), .ck(clk), .q(\cache_data[6][96] )
         );
  dp_1 \cache_data_reg[7][0]  ( .ip(n5935), .ck(clk), .q(\cache_data[7][0] )
         );
  dp_1 \cache_data_reg[7][32]  ( .ip(n5903), .ck(clk), .q(\cache_data[7][32] )
         );
  dp_1 \cache_data_reg[7][64]  ( .ip(n5871), .ck(clk), .q(\cache_data[7][64] )
         );
  dp_1 \cache_data_reg[7][96]  ( .ip(n5839), .ck(clk), .q(\cache_data[7][96] )
         );
  dp_1 \cache_data_reg[8][0]  ( .ip(n5807), .ck(clk), .q(\cache_data[8][0] )
         );
  dp_1 \cache_data_reg[8][32]  ( .ip(n5775), .ck(clk), .q(\cache_data[8][32] )
         );
  dp_1 \cache_data_reg[8][64]  ( .ip(n5743), .ck(clk), .q(\cache_data[8][64] )
         );
  dp_1 \cache_data_reg[8][96]  ( .ip(n5711), .ck(clk), .q(\cache_data[8][96] )
         );
  dp_1 \cache_data_reg[9][0]  ( .ip(n5679), .ck(clk), .q(\cache_data[9][0] )
         );
  dp_1 \cache_data_reg[9][32]  ( .ip(n5647), .ck(clk), .q(\cache_data[9][32] )
         );
  dp_1 \cache_data_reg[9][64]  ( .ip(n5615), .ck(clk), .q(\cache_data[9][64] )
         );
  dp_1 \cache_data_reg[9][96]  ( .ip(n5583), .ck(clk), .q(\cache_data[9][96] )
         );
  dp_1 \cache_data_reg[10][0]  ( .ip(n5551), .ck(clk), .q(\cache_data[10][0] )
         );
  dp_1 \cache_data_reg[10][32]  ( .ip(n5519), .ck(clk), .q(
        \cache_data[10][32] ) );
  dp_1 \cache_data_reg[10][64]  ( .ip(n5487), .ck(clk), .q(
        \cache_data[10][64] ) );
  dp_1 \cache_data_reg[10][96]  ( .ip(n5455), .ck(clk), .q(
        \cache_data[10][96] ) );
  dp_1 \cache_data_reg[11][0]  ( .ip(n5423), .ck(clk), .q(\cache_data[11][0] )
         );
  dp_1 \cache_data_reg[11][32]  ( .ip(n5391), .ck(clk), .q(
        \cache_data[11][32] ) );
  dp_1 \cache_data_reg[11][64]  ( .ip(n5359), .ck(clk), .q(
        \cache_data[11][64] ) );
  dp_1 \cache_data_reg[11][96]  ( .ip(n5327), .ck(clk), .q(
        \cache_data[11][96] ) );
  dp_1 \cache_data_reg[12][0]  ( .ip(n5295), .ck(clk), .q(\cache_data[12][0] )
         );
  dp_1 \cache_data_reg[12][32]  ( .ip(n5263), .ck(clk), .q(
        \cache_data[12][32] ) );
  dp_1 \cache_data_reg[12][64]  ( .ip(n5231), .ck(clk), .q(
        \cache_data[12][64] ) );
  dp_1 \cache_data_reg[12][96]  ( .ip(n5199), .ck(clk), .q(
        \cache_data[12][96] ) );
  dp_1 \cache_data_reg[13][0]  ( .ip(n5167), .ck(clk), .q(\cache_data[13][0] )
         );
  dp_1 \cache_data_reg[13][32]  ( .ip(n5135), .ck(clk), .q(
        \cache_data[13][32] ) );
  dp_1 \cache_data_reg[13][64]  ( .ip(n5103), .ck(clk), .q(
        \cache_data[13][64] ) );
  dp_1 \cache_data_reg[13][96]  ( .ip(n5071), .ck(clk), .q(
        \cache_data[13][96] ) );
  dp_1 \cache_data_reg[14][0]  ( .ip(n5039), .ck(clk), .q(\cache_data[14][0] )
         );
  dp_1 \cache_data_reg[14][32]  ( .ip(n5007), .ck(clk), .q(
        \cache_data[14][32] ) );
  dp_1 \cache_data_reg[14][64]  ( .ip(n4975), .ck(clk), .q(
        \cache_data[14][64] ) );
  dp_1 \cache_data_reg[14][96]  ( .ip(n4943), .ck(clk), .q(
        \cache_data[14][96] ) );
  dp_1 \cache_data_reg[15][0]  ( .ip(n4911), .ck(clk), .q(\cache_data[15][0] )
         );
  dp_1 \cache_data_reg[15][32]  ( .ip(n4879), .ck(clk), .q(
        \cache_data[15][32] ) );
  dp_1 \cache_data_reg[15][64]  ( .ip(n4847), .ck(clk), .q(
        \cache_data[15][64] ) );
  dp_1 \cache_data_reg[15][96]  ( .ip(n4815), .ck(clk), .q(
        \cache_data[15][96] ) );
  dp_1 \iCache_data_wr_reg[1]  ( .ip(n6862), .ck(clk), .q(iCache_data_wr[1])
         );
  dp_1 \cache_data_reg[0][1]  ( .ip(n6830), .ck(clk), .q(\cache_data[0][1] )
         );
  dp_1 \cache_data_reg[0][33]  ( .ip(n6798), .ck(clk), .q(\cache_data[0][33] )
         );
  dp_1 \cache_data_reg[0][65]  ( .ip(n6766), .ck(clk), .q(\cache_data[0][65] )
         );
  dp_1 \cache_data_reg[0][97]  ( .ip(n6734), .ck(clk), .q(\cache_data[0][97] )
         );
  dp_1 \cache_data_reg[1][1]  ( .ip(n6702), .ck(clk), .q(\cache_data[1][1] )
         );
  dp_1 \cache_data_reg[1][33]  ( .ip(n6670), .ck(clk), .q(\cache_data[1][33] )
         );
  dp_1 \cache_data_reg[1][65]  ( .ip(n6638), .ck(clk), .q(\cache_data[1][65] )
         );
  dp_1 \cache_data_reg[1][97]  ( .ip(n6606), .ck(clk), .q(\cache_data[1][97] )
         );
  dp_1 \cache_data_reg[2][1]  ( .ip(n6574), .ck(clk), .q(\cache_data[2][1] )
         );
  dp_1 \cache_data_reg[2][33]  ( .ip(n6542), .ck(clk), .q(\cache_data[2][33] )
         );
  dp_1 \cache_data_reg[2][65]  ( .ip(n6510), .ck(clk), .q(\cache_data[2][65] )
         );
  dp_1 \cache_data_reg[2][97]  ( .ip(n6478), .ck(clk), .q(\cache_data[2][97] )
         );
  dp_1 \cache_data_reg[3][1]  ( .ip(n6446), .ck(clk), .q(\cache_data[3][1] )
         );
  dp_1 \cache_data_reg[3][33]  ( .ip(n6414), .ck(clk), .q(\cache_data[3][33] )
         );
  dp_1 \cache_data_reg[3][65]  ( .ip(n6382), .ck(clk), .q(\cache_data[3][65] )
         );
  dp_1 \cache_data_reg[3][97]  ( .ip(n6350), .ck(clk), .q(\cache_data[3][97] )
         );
  dp_1 \cache_data_reg[4][1]  ( .ip(n6318), .ck(clk), .q(\cache_data[4][1] )
         );
  dp_1 \cache_data_reg[4][33]  ( .ip(n6286), .ck(clk), .q(\cache_data[4][33] )
         );
  dp_1 \cache_data_reg[4][65]  ( .ip(n6254), .ck(clk), .q(\cache_data[4][65] )
         );
  dp_1 \cache_data_reg[4][97]  ( .ip(n6222), .ck(clk), .q(\cache_data[4][97] )
         );
  dp_1 \cache_data_reg[5][1]  ( .ip(n6190), .ck(clk), .q(\cache_data[5][1] )
         );
  dp_1 \cache_data_reg[5][33]  ( .ip(n6158), .ck(clk), .q(\cache_data[5][33] )
         );
  dp_1 \cache_data_reg[5][65]  ( .ip(n6126), .ck(clk), .q(\cache_data[5][65] )
         );
  dp_1 \cache_data_reg[5][97]  ( .ip(n6094), .ck(clk), .q(\cache_data[5][97] )
         );
  dp_1 \cache_data_reg[6][1]  ( .ip(n6062), .ck(clk), .q(\cache_data[6][1] )
         );
  dp_1 \cache_data_reg[6][33]  ( .ip(n6030), .ck(clk), .q(\cache_data[6][33] )
         );
  dp_1 \cache_data_reg[6][65]  ( .ip(n5998), .ck(clk), .q(\cache_data[6][65] )
         );
  dp_1 \cache_data_reg[6][97]  ( .ip(n5966), .ck(clk), .q(\cache_data[6][97] )
         );
  dp_1 \cache_data_reg[7][1]  ( .ip(n5934), .ck(clk), .q(\cache_data[7][1] )
         );
  dp_1 \cache_data_reg[7][33]  ( .ip(n5902), .ck(clk), .q(\cache_data[7][33] )
         );
  dp_1 \cache_data_reg[7][65]  ( .ip(n5870), .ck(clk), .q(\cache_data[7][65] )
         );
  dp_1 \cache_data_reg[7][97]  ( .ip(n5838), .ck(clk), .q(\cache_data[7][97] )
         );
  dp_1 \cache_data_reg[8][1]  ( .ip(n5806), .ck(clk), .q(\cache_data[8][1] )
         );
  dp_1 \cache_data_reg[8][33]  ( .ip(n5774), .ck(clk), .q(\cache_data[8][33] )
         );
  dp_1 \cache_data_reg[8][65]  ( .ip(n5742), .ck(clk), .q(\cache_data[8][65] )
         );
  dp_1 \cache_data_reg[8][97]  ( .ip(n5710), .ck(clk), .q(\cache_data[8][97] )
         );
  dp_1 \cache_data_reg[9][1]  ( .ip(n5678), .ck(clk), .q(\cache_data[9][1] )
         );
  dp_1 \cache_data_reg[9][33]  ( .ip(n5646), .ck(clk), .q(\cache_data[9][33] )
         );
  dp_1 \cache_data_reg[9][65]  ( .ip(n5614), .ck(clk), .q(\cache_data[9][65] )
         );
  dp_1 \cache_data_reg[9][97]  ( .ip(n5582), .ck(clk), .q(\cache_data[9][97] )
         );
  dp_1 \cache_data_reg[10][1]  ( .ip(n5550), .ck(clk), .q(\cache_data[10][1] )
         );
  dp_1 \cache_data_reg[10][33]  ( .ip(n5518), .ck(clk), .q(
        \cache_data[10][33] ) );
  dp_1 \cache_data_reg[10][65]  ( .ip(n5486), .ck(clk), .q(
        \cache_data[10][65] ) );
  dp_1 \cache_data_reg[10][97]  ( .ip(n5454), .ck(clk), .q(
        \cache_data[10][97] ) );
  dp_1 \cache_data_reg[11][1]  ( .ip(n5422), .ck(clk), .q(\cache_data[11][1] )
         );
  dp_1 \cache_data_reg[11][33]  ( .ip(n5390), .ck(clk), .q(
        \cache_data[11][33] ) );
  dp_1 \cache_data_reg[11][65]  ( .ip(n5358), .ck(clk), .q(
        \cache_data[11][65] ) );
  dp_1 \cache_data_reg[11][97]  ( .ip(n5326), .ck(clk), .q(
        \cache_data[11][97] ) );
  dp_1 \cache_data_reg[12][1]  ( .ip(n5294), .ck(clk), .q(\cache_data[12][1] )
         );
  dp_1 \cache_data_reg[12][33]  ( .ip(n5262), .ck(clk), .q(
        \cache_data[12][33] ) );
  dp_1 \cache_data_reg[12][65]  ( .ip(n5230), .ck(clk), .q(
        \cache_data[12][65] ) );
  dp_1 \cache_data_reg[12][97]  ( .ip(n5198), .ck(clk), .q(
        \cache_data[12][97] ) );
  dp_1 \cache_data_reg[13][1]  ( .ip(n5166), .ck(clk), .q(\cache_data[13][1] )
         );
  dp_1 \cache_data_reg[13][33]  ( .ip(n5134), .ck(clk), .q(
        \cache_data[13][33] ) );
  dp_1 \cache_data_reg[13][65]  ( .ip(n5102), .ck(clk), .q(
        \cache_data[13][65] ) );
  dp_1 \cache_data_reg[13][97]  ( .ip(n5070), .ck(clk), .q(
        \cache_data[13][97] ) );
  dp_1 \cache_data_reg[14][1]  ( .ip(n5038), .ck(clk), .q(\cache_data[14][1] )
         );
  dp_1 \cache_data_reg[14][33]  ( .ip(n5006), .ck(clk), .q(
        \cache_data[14][33] ) );
  dp_1 \cache_data_reg[14][65]  ( .ip(n4974), .ck(clk), .q(
        \cache_data[14][65] ) );
  dp_1 \cache_data_reg[14][97]  ( .ip(n4942), .ck(clk), .q(
        \cache_data[14][97] ) );
  dp_1 \cache_data_reg[15][1]  ( .ip(n4910), .ck(clk), .q(\cache_data[15][1] )
         );
  dp_1 \cache_data_reg[15][33]  ( .ip(n4878), .ck(clk), .q(
        \cache_data[15][33] ) );
  dp_1 \cache_data_reg[15][65]  ( .ip(n4846), .ck(clk), .q(
        \cache_data[15][65] ) );
  dp_1 \cache_data_reg[15][97]  ( .ip(n4814), .ck(clk), .q(
        \cache_data[15][97] ) );
  dp_1 \iCache_data_wr_reg[2]  ( .ip(n6861), .ck(clk), .q(iCache_data_wr[2])
         );
  dp_1 \cache_data_reg[0][2]  ( .ip(n6829), .ck(clk), .q(\cache_data[0][2] )
         );
  dp_1 \cache_data_reg[0][34]  ( .ip(n6797), .ck(clk), .q(\cache_data[0][34] )
         );
  dp_1 \cache_data_reg[0][66]  ( .ip(n6765), .ck(clk), .q(\cache_data[0][66] )
         );
  dp_1 \cache_data_reg[0][98]  ( .ip(n6733), .ck(clk), .q(\cache_data[0][98] )
         );
  dp_1 \cache_data_reg[1][2]  ( .ip(n6701), .ck(clk), .q(\cache_data[1][2] )
         );
  dp_1 \cache_data_reg[1][34]  ( .ip(n6669), .ck(clk), .q(\cache_data[1][34] )
         );
  dp_1 \cache_data_reg[1][66]  ( .ip(n6637), .ck(clk), .q(\cache_data[1][66] )
         );
  dp_1 \cache_data_reg[1][98]  ( .ip(n6605), .ck(clk), .q(\cache_data[1][98] )
         );
  dp_1 \cache_data_reg[2][2]  ( .ip(n6573), .ck(clk), .q(\cache_data[2][2] )
         );
  dp_1 \cache_data_reg[2][34]  ( .ip(n6541), .ck(clk), .q(\cache_data[2][34] )
         );
  dp_1 \cache_data_reg[2][66]  ( .ip(n6509), .ck(clk), .q(\cache_data[2][66] )
         );
  dp_1 \cache_data_reg[2][98]  ( .ip(n6477), .ck(clk), .q(\cache_data[2][98] )
         );
  dp_1 \cache_data_reg[3][2]  ( .ip(n6445), .ck(clk), .q(\cache_data[3][2] )
         );
  dp_1 \cache_data_reg[3][34]  ( .ip(n6413), .ck(clk), .q(\cache_data[3][34] )
         );
  dp_1 \cache_data_reg[3][66]  ( .ip(n6381), .ck(clk), .q(\cache_data[3][66] )
         );
  dp_1 \cache_data_reg[3][98]  ( .ip(n6349), .ck(clk), .q(\cache_data[3][98] )
         );
  dp_1 \cache_data_reg[4][2]  ( .ip(n6317), .ck(clk), .q(\cache_data[4][2] )
         );
  dp_1 \cache_data_reg[4][34]  ( .ip(n6285), .ck(clk), .q(\cache_data[4][34] )
         );
  dp_1 \cache_data_reg[4][66]  ( .ip(n6253), .ck(clk), .q(\cache_data[4][66] )
         );
  dp_1 \cache_data_reg[4][98]  ( .ip(n6221), .ck(clk), .q(\cache_data[4][98] )
         );
  dp_1 \cache_data_reg[5][2]  ( .ip(n6189), .ck(clk), .q(\cache_data[5][2] )
         );
  dp_1 \cache_data_reg[5][34]  ( .ip(n6157), .ck(clk), .q(\cache_data[5][34] )
         );
  dp_1 \cache_data_reg[5][66]  ( .ip(n6125), .ck(clk), .q(\cache_data[5][66] )
         );
  dp_1 \cache_data_reg[5][98]  ( .ip(n6093), .ck(clk), .q(\cache_data[5][98] )
         );
  dp_1 \cache_data_reg[6][2]  ( .ip(n6061), .ck(clk), .q(\cache_data[6][2] )
         );
  dp_1 \cache_data_reg[6][34]  ( .ip(n6029), .ck(clk), .q(\cache_data[6][34] )
         );
  dp_1 \cache_data_reg[6][66]  ( .ip(n5997), .ck(clk), .q(\cache_data[6][66] )
         );
  dp_1 \cache_data_reg[6][98]  ( .ip(n5965), .ck(clk), .q(\cache_data[6][98] )
         );
  dp_1 \cache_data_reg[7][2]  ( .ip(n5933), .ck(clk), .q(\cache_data[7][2] )
         );
  dp_1 \cache_data_reg[7][34]  ( .ip(n5901), .ck(clk), .q(\cache_data[7][34] )
         );
  dp_1 \cache_data_reg[7][66]  ( .ip(n5869), .ck(clk), .q(\cache_data[7][66] )
         );
  dp_1 \cache_data_reg[7][98]  ( .ip(n5837), .ck(clk), .q(\cache_data[7][98] )
         );
  dp_1 \cache_data_reg[8][2]  ( .ip(n5805), .ck(clk), .q(\cache_data[8][2] )
         );
  dp_1 \cache_data_reg[8][34]  ( .ip(n5773), .ck(clk), .q(\cache_data[8][34] )
         );
  dp_1 \cache_data_reg[8][66]  ( .ip(n5741), .ck(clk), .q(\cache_data[8][66] )
         );
  dp_1 \cache_data_reg[8][98]  ( .ip(n5709), .ck(clk), .q(\cache_data[8][98] )
         );
  dp_1 \cache_data_reg[9][2]  ( .ip(n5677), .ck(clk), .q(\cache_data[9][2] )
         );
  dp_1 \cache_data_reg[9][34]  ( .ip(n5645), .ck(clk), .q(\cache_data[9][34] )
         );
  dp_1 \cache_data_reg[9][66]  ( .ip(n5613), .ck(clk), .q(\cache_data[9][66] )
         );
  dp_1 \cache_data_reg[9][98]  ( .ip(n5581), .ck(clk), .q(\cache_data[9][98] )
         );
  dp_1 \cache_data_reg[10][2]  ( .ip(n5549), .ck(clk), .q(\cache_data[10][2] )
         );
  dp_1 \cache_data_reg[10][34]  ( .ip(n5517), .ck(clk), .q(
        \cache_data[10][34] ) );
  dp_1 \cache_data_reg[10][66]  ( .ip(n5485), .ck(clk), .q(
        \cache_data[10][66] ) );
  dp_1 \cache_data_reg[10][98]  ( .ip(n5453), .ck(clk), .q(
        \cache_data[10][98] ) );
  dp_1 \cache_data_reg[11][2]  ( .ip(n5421), .ck(clk), .q(\cache_data[11][2] )
         );
  dp_1 \cache_data_reg[11][34]  ( .ip(n5389), .ck(clk), .q(
        \cache_data[11][34] ) );
  dp_1 \cache_data_reg[11][66]  ( .ip(n5357), .ck(clk), .q(
        \cache_data[11][66] ) );
  dp_1 \cache_data_reg[11][98]  ( .ip(n5325), .ck(clk), .q(
        \cache_data[11][98] ) );
  dp_1 \cache_data_reg[12][2]  ( .ip(n5293), .ck(clk), .q(\cache_data[12][2] )
         );
  dp_1 \cache_data_reg[12][34]  ( .ip(n5261), .ck(clk), .q(
        \cache_data[12][34] ) );
  dp_1 \cache_data_reg[12][66]  ( .ip(n5229), .ck(clk), .q(
        \cache_data[12][66] ) );
  dp_1 \cache_data_reg[12][98]  ( .ip(n5197), .ck(clk), .q(
        \cache_data[12][98] ) );
  dp_1 \cache_data_reg[13][2]  ( .ip(n5165), .ck(clk), .q(\cache_data[13][2] )
         );
  dp_1 \cache_data_reg[13][34]  ( .ip(n5133), .ck(clk), .q(
        \cache_data[13][34] ) );
  dp_1 \cache_data_reg[13][66]  ( .ip(n5101), .ck(clk), .q(
        \cache_data[13][66] ) );
  dp_1 \cache_data_reg[13][98]  ( .ip(n5069), .ck(clk), .q(
        \cache_data[13][98] ) );
  dp_1 \cache_data_reg[14][2]  ( .ip(n5037), .ck(clk), .q(\cache_data[14][2] )
         );
  dp_1 \cache_data_reg[14][34]  ( .ip(n5005), .ck(clk), .q(
        \cache_data[14][34] ) );
  dp_1 \cache_data_reg[14][66]  ( .ip(n4973), .ck(clk), .q(
        \cache_data[14][66] ) );
  dp_1 \cache_data_reg[14][98]  ( .ip(n4941), .ck(clk), .q(
        \cache_data[14][98] ) );
  dp_1 \cache_data_reg[15][2]  ( .ip(n4909), .ck(clk), .q(\cache_data[15][2] )
         );
  dp_1 \cache_data_reg[15][34]  ( .ip(n4877), .ck(clk), .q(
        \cache_data[15][34] ) );
  dp_1 \cache_data_reg[15][66]  ( .ip(n4845), .ck(clk), .q(
        \cache_data[15][66] ) );
  dp_1 \cache_data_reg[15][98]  ( .ip(n4813), .ck(clk), .q(
        \cache_data[15][98] ) );
  dp_1 \iCache_data_wr_reg[3]  ( .ip(n6860), .ck(clk), .q(iCache_data_wr[3])
         );
  dp_1 \cache_data_reg[0][3]  ( .ip(n6828), .ck(clk), .q(\cache_data[0][3] )
         );
  dp_1 \cache_data_reg[0][35]  ( .ip(n6796), .ck(clk), .q(\cache_data[0][35] )
         );
  dp_1 \cache_data_reg[0][67]  ( .ip(n6764), .ck(clk), .q(\cache_data[0][67] )
         );
  dp_1 \cache_data_reg[0][99]  ( .ip(n6732), .ck(clk), .q(\cache_data[0][99] )
         );
  dp_1 \cache_data_reg[1][3]  ( .ip(n6700), .ck(clk), .q(\cache_data[1][3] )
         );
  dp_1 \cache_data_reg[1][35]  ( .ip(n6668), .ck(clk), .q(\cache_data[1][35] )
         );
  dp_1 \cache_data_reg[1][67]  ( .ip(n6636), .ck(clk), .q(\cache_data[1][67] )
         );
  dp_1 \cache_data_reg[1][99]  ( .ip(n6604), .ck(clk), .q(\cache_data[1][99] )
         );
  dp_1 \cache_data_reg[2][3]  ( .ip(n6572), .ck(clk), .q(\cache_data[2][3] )
         );
  dp_1 \cache_data_reg[2][35]  ( .ip(n6540), .ck(clk), .q(\cache_data[2][35] )
         );
  dp_1 \cache_data_reg[2][67]  ( .ip(n6508), .ck(clk), .q(\cache_data[2][67] )
         );
  dp_1 \cache_data_reg[2][99]  ( .ip(n6476), .ck(clk), .q(\cache_data[2][99] )
         );
  dp_1 \cache_data_reg[3][3]  ( .ip(n6444), .ck(clk), .q(\cache_data[3][3] )
         );
  dp_1 \cache_data_reg[3][35]  ( .ip(n6412), .ck(clk), .q(\cache_data[3][35] )
         );
  dp_1 \cache_data_reg[3][67]  ( .ip(n6380), .ck(clk), .q(\cache_data[3][67] )
         );
  dp_1 \cache_data_reg[3][99]  ( .ip(n6348), .ck(clk), .q(\cache_data[3][99] )
         );
  dp_1 \cache_data_reg[4][3]  ( .ip(n6316), .ck(clk), .q(\cache_data[4][3] )
         );
  dp_1 \cache_data_reg[4][35]  ( .ip(n6284), .ck(clk), .q(\cache_data[4][35] )
         );
  dp_1 \cache_data_reg[4][67]  ( .ip(n6252), .ck(clk), .q(\cache_data[4][67] )
         );
  dp_1 \cache_data_reg[4][99]  ( .ip(n6220), .ck(clk), .q(\cache_data[4][99] )
         );
  dp_1 \cache_data_reg[5][3]  ( .ip(n6188), .ck(clk), .q(\cache_data[5][3] )
         );
  dp_1 \cache_data_reg[5][35]  ( .ip(n6156), .ck(clk), .q(\cache_data[5][35] )
         );
  dp_1 \cache_data_reg[5][67]  ( .ip(n6124), .ck(clk), .q(\cache_data[5][67] )
         );
  dp_1 \cache_data_reg[5][99]  ( .ip(n6092), .ck(clk), .q(\cache_data[5][99] )
         );
  dp_1 \cache_data_reg[6][3]  ( .ip(n6060), .ck(clk), .q(\cache_data[6][3] )
         );
  dp_1 \cache_data_reg[6][35]  ( .ip(n6028), .ck(clk), .q(\cache_data[6][35] )
         );
  dp_1 \cache_data_reg[6][67]  ( .ip(n5996), .ck(clk), .q(\cache_data[6][67] )
         );
  dp_1 \cache_data_reg[6][99]  ( .ip(n5964), .ck(clk), .q(\cache_data[6][99] )
         );
  dp_1 \cache_data_reg[7][3]  ( .ip(n5932), .ck(clk), .q(\cache_data[7][3] )
         );
  dp_1 \cache_data_reg[7][35]  ( .ip(n5900), .ck(clk), .q(\cache_data[7][35] )
         );
  dp_1 \cache_data_reg[7][67]  ( .ip(n5868), .ck(clk), .q(\cache_data[7][67] )
         );
  dp_1 \cache_data_reg[7][99]  ( .ip(n5836), .ck(clk), .q(\cache_data[7][99] )
         );
  dp_1 \cache_data_reg[8][3]  ( .ip(n5804), .ck(clk), .q(\cache_data[8][3] )
         );
  dp_1 \cache_data_reg[8][35]  ( .ip(n5772), .ck(clk), .q(\cache_data[8][35] )
         );
  dp_1 \cache_data_reg[8][67]  ( .ip(n5740), .ck(clk), .q(\cache_data[8][67] )
         );
  dp_1 \cache_data_reg[8][99]  ( .ip(n5708), .ck(clk), .q(\cache_data[8][99] )
         );
  dp_1 \cache_data_reg[9][3]  ( .ip(n5676), .ck(clk), .q(\cache_data[9][3] )
         );
  dp_1 \cache_data_reg[9][35]  ( .ip(n5644), .ck(clk), .q(\cache_data[9][35] )
         );
  dp_1 \cache_data_reg[9][67]  ( .ip(n5612), .ck(clk), .q(\cache_data[9][67] )
         );
  dp_1 \cache_data_reg[9][99]  ( .ip(n5580), .ck(clk), .q(\cache_data[9][99] )
         );
  dp_1 \cache_data_reg[10][3]  ( .ip(n5548), .ck(clk), .q(\cache_data[10][3] )
         );
  dp_1 \cache_data_reg[10][35]  ( .ip(n5516), .ck(clk), .q(
        \cache_data[10][35] ) );
  dp_1 \cache_data_reg[10][67]  ( .ip(n5484), .ck(clk), .q(
        \cache_data[10][67] ) );
  dp_1 \cache_data_reg[10][99]  ( .ip(n5452), .ck(clk), .q(
        \cache_data[10][99] ) );
  dp_1 \cache_data_reg[11][3]  ( .ip(n5420), .ck(clk), .q(\cache_data[11][3] )
         );
  dp_1 \cache_data_reg[11][35]  ( .ip(n5388), .ck(clk), .q(
        \cache_data[11][35] ) );
  dp_1 \cache_data_reg[11][67]  ( .ip(n5356), .ck(clk), .q(
        \cache_data[11][67] ) );
  dp_1 \cache_data_reg[11][99]  ( .ip(n5324), .ck(clk), .q(
        \cache_data[11][99] ) );
  dp_1 \cache_data_reg[12][3]  ( .ip(n5292), .ck(clk), .q(\cache_data[12][3] )
         );
  dp_1 \cache_data_reg[12][35]  ( .ip(n5260), .ck(clk), .q(
        \cache_data[12][35] ) );
  dp_1 \cache_data_reg[12][67]  ( .ip(n5228), .ck(clk), .q(
        \cache_data[12][67] ) );
  dp_1 \cache_data_reg[12][99]  ( .ip(n5196), .ck(clk), .q(
        \cache_data[12][99] ) );
  dp_1 \cache_data_reg[13][3]  ( .ip(n5164), .ck(clk), .q(\cache_data[13][3] )
         );
  dp_1 \cache_data_reg[13][35]  ( .ip(n5132), .ck(clk), .q(
        \cache_data[13][35] ) );
  dp_1 \cache_data_reg[13][67]  ( .ip(n5100), .ck(clk), .q(
        \cache_data[13][67] ) );
  dp_1 \cache_data_reg[13][99]  ( .ip(n5068), .ck(clk), .q(
        \cache_data[13][99] ) );
  dp_1 \cache_data_reg[14][3]  ( .ip(n5036), .ck(clk), .q(\cache_data[14][3] )
         );
  dp_1 \cache_data_reg[14][35]  ( .ip(n5004), .ck(clk), .q(
        \cache_data[14][35] ) );
  dp_1 \cache_data_reg[14][67]  ( .ip(n4972), .ck(clk), .q(
        \cache_data[14][67] ) );
  dp_1 \cache_data_reg[14][99]  ( .ip(n4940), .ck(clk), .q(
        \cache_data[14][99] ) );
  dp_1 \cache_data_reg[15][3]  ( .ip(n4908), .ck(clk), .q(\cache_data[15][3] )
         );
  dp_1 \cache_data_reg[15][35]  ( .ip(n4876), .ck(clk), .q(
        \cache_data[15][35] ) );
  dp_1 \cache_data_reg[15][67]  ( .ip(n4844), .ck(clk), .q(
        \cache_data[15][67] ) );
  dp_1 \cache_data_reg[15][99]  ( .ip(n4812), .ck(clk), .q(
        \cache_data[15][99] ) );
  dp_1 \iCache_data_wr_reg[4]  ( .ip(n6859), .ck(clk), .q(iCache_data_wr[4])
         );
  dp_1 \cache_data_reg[0][4]  ( .ip(n6827), .ck(clk), .q(\cache_data[0][4] )
         );
  dp_1 \cache_data_reg[0][36]  ( .ip(n6795), .ck(clk), .q(\cache_data[0][36] )
         );
  dp_1 \cache_data_reg[0][68]  ( .ip(n6763), .ck(clk), .q(\cache_data[0][68] )
         );
  dp_1 \cache_data_reg[0][100]  ( .ip(n6731), .ck(clk), .q(
        \cache_data[0][100] ) );
  dp_1 \cache_data_reg[1][4]  ( .ip(n6699), .ck(clk), .q(\cache_data[1][4] )
         );
  dp_1 \cache_data_reg[1][36]  ( .ip(n6667), .ck(clk), .q(\cache_data[1][36] )
         );
  dp_1 \cache_data_reg[1][68]  ( .ip(n6635), .ck(clk), .q(\cache_data[1][68] )
         );
  dp_1 \cache_data_reg[1][100]  ( .ip(n6603), .ck(clk), .q(
        \cache_data[1][100] ) );
  dp_1 \cache_data_reg[2][4]  ( .ip(n6571), .ck(clk), .q(\cache_data[2][4] )
         );
  dp_1 \cache_data_reg[2][36]  ( .ip(n6539), .ck(clk), .q(\cache_data[2][36] )
         );
  dp_1 \cache_data_reg[2][68]  ( .ip(n6507), .ck(clk), .q(\cache_data[2][68] )
         );
  dp_1 \cache_data_reg[2][100]  ( .ip(n6475), .ck(clk), .q(
        \cache_data[2][100] ) );
  dp_1 \cache_data_reg[3][4]  ( .ip(n6443), .ck(clk), .q(\cache_data[3][4] )
         );
  dp_1 \cache_data_reg[3][36]  ( .ip(n6411), .ck(clk), .q(\cache_data[3][36] )
         );
  dp_1 \cache_data_reg[3][68]  ( .ip(n6379), .ck(clk), .q(\cache_data[3][68] )
         );
  dp_1 \cache_data_reg[3][100]  ( .ip(n6347), .ck(clk), .q(
        \cache_data[3][100] ) );
  dp_1 \cache_data_reg[4][4]  ( .ip(n6315), .ck(clk), .q(\cache_data[4][4] )
         );
  dp_1 \cache_data_reg[4][36]  ( .ip(n6283), .ck(clk), .q(\cache_data[4][36] )
         );
  dp_1 \cache_data_reg[4][68]  ( .ip(n6251), .ck(clk), .q(\cache_data[4][68] )
         );
  dp_1 \cache_data_reg[4][100]  ( .ip(n6219), .ck(clk), .q(
        \cache_data[4][100] ) );
  dp_1 \cache_data_reg[5][4]  ( .ip(n6187), .ck(clk), .q(\cache_data[5][4] )
         );
  dp_1 \cache_data_reg[5][36]  ( .ip(n6155), .ck(clk), .q(\cache_data[5][36] )
         );
  dp_1 \cache_data_reg[5][68]  ( .ip(n6123), .ck(clk), .q(\cache_data[5][68] )
         );
  dp_1 \cache_data_reg[5][100]  ( .ip(n6091), .ck(clk), .q(
        \cache_data[5][100] ) );
  dp_1 \cache_data_reg[6][4]  ( .ip(n6059), .ck(clk), .q(\cache_data[6][4] )
         );
  dp_1 \cache_data_reg[6][36]  ( .ip(n6027), .ck(clk), .q(\cache_data[6][36] )
         );
  dp_1 \cache_data_reg[6][68]  ( .ip(n5995), .ck(clk), .q(\cache_data[6][68] )
         );
  dp_1 \cache_data_reg[6][100]  ( .ip(n5963), .ck(clk), .q(
        \cache_data[6][100] ) );
  dp_1 \cache_data_reg[7][4]  ( .ip(n5931), .ck(clk), .q(\cache_data[7][4] )
         );
  dp_1 \cache_data_reg[7][36]  ( .ip(n5899), .ck(clk), .q(\cache_data[7][36] )
         );
  dp_1 \cache_data_reg[7][68]  ( .ip(n5867), .ck(clk), .q(\cache_data[7][68] )
         );
  dp_1 \cache_data_reg[7][100]  ( .ip(n5835), .ck(clk), .q(
        \cache_data[7][100] ) );
  dp_1 \cache_data_reg[8][4]  ( .ip(n5803), .ck(clk), .q(\cache_data[8][4] )
         );
  dp_1 \cache_data_reg[8][36]  ( .ip(n5771), .ck(clk), .q(\cache_data[8][36] )
         );
  dp_1 \cache_data_reg[8][68]  ( .ip(n5739), .ck(clk), .q(\cache_data[8][68] )
         );
  dp_1 \cache_data_reg[8][100]  ( .ip(n5707), .ck(clk), .q(
        \cache_data[8][100] ) );
  dp_1 \cache_data_reg[9][4]  ( .ip(n5675), .ck(clk), .q(\cache_data[9][4] )
         );
  dp_1 \cache_data_reg[9][36]  ( .ip(n5643), .ck(clk), .q(\cache_data[9][36] )
         );
  dp_1 \cache_data_reg[9][68]  ( .ip(n5611), .ck(clk), .q(\cache_data[9][68] )
         );
  dp_1 \cache_data_reg[9][100]  ( .ip(n5579), .ck(clk), .q(
        \cache_data[9][100] ) );
  dp_1 \cache_data_reg[10][4]  ( .ip(n5547), .ck(clk), .q(\cache_data[10][4] )
         );
  dp_1 \cache_data_reg[10][36]  ( .ip(n5515), .ck(clk), .q(
        \cache_data[10][36] ) );
  dp_1 \cache_data_reg[10][68]  ( .ip(n5483), .ck(clk), .q(
        \cache_data[10][68] ) );
  dp_1 \cache_data_reg[10][100]  ( .ip(n5451), .ck(clk), .q(
        \cache_data[10][100] ) );
  dp_1 \cache_data_reg[11][4]  ( .ip(n5419), .ck(clk), .q(\cache_data[11][4] )
         );
  dp_1 \cache_data_reg[11][36]  ( .ip(n5387), .ck(clk), .q(
        \cache_data[11][36] ) );
  dp_1 \cache_data_reg[11][68]  ( .ip(n5355), .ck(clk), .q(
        \cache_data[11][68] ) );
  dp_1 \cache_data_reg[11][100]  ( .ip(n5323), .ck(clk), .q(
        \cache_data[11][100] ) );
  dp_1 \cache_data_reg[12][4]  ( .ip(n5291), .ck(clk), .q(\cache_data[12][4] )
         );
  dp_1 \cache_data_reg[12][36]  ( .ip(n5259), .ck(clk), .q(
        \cache_data[12][36] ) );
  dp_1 \cache_data_reg[12][68]  ( .ip(n5227), .ck(clk), .q(
        \cache_data[12][68] ) );
  dp_1 \cache_data_reg[12][100]  ( .ip(n5195), .ck(clk), .q(
        \cache_data[12][100] ) );
  dp_1 \cache_data_reg[13][4]  ( .ip(n5163), .ck(clk), .q(\cache_data[13][4] )
         );
  dp_1 \cache_data_reg[13][36]  ( .ip(n5131), .ck(clk), .q(
        \cache_data[13][36] ) );
  dp_1 \cache_data_reg[13][68]  ( .ip(n5099), .ck(clk), .q(
        \cache_data[13][68] ) );
  dp_1 \cache_data_reg[13][100]  ( .ip(n5067), .ck(clk), .q(
        \cache_data[13][100] ) );
  dp_1 \cache_data_reg[14][4]  ( .ip(n5035), .ck(clk), .q(\cache_data[14][4] )
         );
  dp_1 \cache_data_reg[14][36]  ( .ip(n5003), .ck(clk), .q(
        \cache_data[14][36] ) );
  dp_1 \cache_data_reg[14][68]  ( .ip(n4971), .ck(clk), .q(
        \cache_data[14][68] ) );
  dp_1 \cache_data_reg[14][100]  ( .ip(n4939), .ck(clk), .q(
        \cache_data[14][100] ) );
  dp_1 \cache_data_reg[15][4]  ( .ip(n4907), .ck(clk), .q(\cache_data[15][4] )
         );
  dp_1 \cache_data_reg[15][36]  ( .ip(n4875), .ck(clk), .q(
        \cache_data[15][36] ) );
  dp_1 \cache_data_reg[15][68]  ( .ip(n4843), .ck(clk), .q(
        \cache_data[15][68] ) );
  dp_1 \cache_data_reg[15][100]  ( .ip(n4811), .ck(clk), .q(
        \cache_data[15][100] ) );
  dp_1 \iCache_data_wr_reg[5]  ( .ip(n6858), .ck(clk), .q(iCache_data_wr[5])
         );
  dp_1 \cache_data_reg[0][5]  ( .ip(n6826), .ck(clk), .q(\cache_data[0][5] )
         );
  dp_1 \cache_data_reg[0][37]  ( .ip(n6794), .ck(clk), .q(\cache_data[0][37] )
         );
  dp_1 \cache_data_reg[0][69]  ( .ip(n6762), .ck(clk), .q(\cache_data[0][69] )
         );
  dp_1 \cache_data_reg[0][101]  ( .ip(n6730), .ck(clk), .q(
        \cache_data[0][101] ) );
  dp_1 \cache_data_reg[1][5]  ( .ip(n6698), .ck(clk), .q(\cache_data[1][5] )
         );
  dp_1 \cache_data_reg[1][37]  ( .ip(n6666), .ck(clk), .q(\cache_data[1][37] )
         );
  dp_1 \cache_data_reg[1][69]  ( .ip(n6634), .ck(clk), .q(\cache_data[1][69] )
         );
  dp_1 \cache_data_reg[1][101]  ( .ip(n6602), .ck(clk), .q(
        \cache_data[1][101] ) );
  dp_1 \cache_data_reg[2][5]  ( .ip(n6570), .ck(clk), .q(\cache_data[2][5] )
         );
  dp_1 \cache_data_reg[2][37]  ( .ip(n6538), .ck(clk), .q(\cache_data[2][37] )
         );
  dp_1 \cache_data_reg[2][69]  ( .ip(n6506), .ck(clk), .q(\cache_data[2][69] )
         );
  dp_1 \cache_data_reg[2][101]  ( .ip(n6474), .ck(clk), .q(
        \cache_data[2][101] ) );
  dp_1 \cache_data_reg[3][5]  ( .ip(n6442), .ck(clk), .q(\cache_data[3][5] )
         );
  dp_1 \cache_data_reg[3][37]  ( .ip(n6410), .ck(clk), .q(\cache_data[3][37] )
         );
  dp_1 \cache_data_reg[3][69]  ( .ip(n6378), .ck(clk), .q(\cache_data[3][69] )
         );
  dp_1 \cache_data_reg[3][101]  ( .ip(n6346), .ck(clk), .q(
        \cache_data[3][101] ) );
  dp_1 \cache_data_reg[4][5]  ( .ip(n6314), .ck(clk), .q(\cache_data[4][5] )
         );
  dp_1 \cache_data_reg[4][37]  ( .ip(n6282), .ck(clk), .q(\cache_data[4][37] )
         );
  dp_1 \cache_data_reg[4][69]  ( .ip(n6250), .ck(clk), .q(\cache_data[4][69] )
         );
  dp_1 \cache_data_reg[4][101]  ( .ip(n6218), .ck(clk), .q(
        \cache_data[4][101] ) );
  dp_1 \cache_data_reg[5][5]  ( .ip(n6186), .ck(clk), .q(\cache_data[5][5] )
         );
  dp_1 \cache_data_reg[5][37]  ( .ip(n6154), .ck(clk), .q(\cache_data[5][37] )
         );
  dp_1 \cache_data_reg[5][69]  ( .ip(n6122), .ck(clk), .q(\cache_data[5][69] )
         );
  dp_1 \cache_data_reg[5][101]  ( .ip(n6090), .ck(clk), .q(
        \cache_data[5][101] ) );
  dp_1 \cache_data_reg[6][5]  ( .ip(n6058), .ck(clk), .q(\cache_data[6][5] )
         );
  dp_1 \cache_data_reg[6][37]  ( .ip(n6026), .ck(clk), .q(\cache_data[6][37] )
         );
  dp_1 \cache_data_reg[6][69]  ( .ip(n5994), .ck(clk), .q(\cache_data[6][69] )
         );
  dp_1 \cache_data_reg[6][101]  ( .ip(n5962), .ck(clk), .q(
        \cache_data[6][101] ) );
  dp_1 \cache_data_reg[7][5]  ( .ip(n5930), .ck(clk), .q(\cache_data[7][5] )
         );
  dp_1 \cache_data_reg[7][37]  ( .ip(n5898), .ck(clk), .q(\cache_data[7][37] )
         );
  dp_1 \cache_data_reg[7][69]  ( .ip(n5866), .ck(clk), .q(\cache_data[7][69] )
         );
  dp_1 \cache_data_reg[7][101]  ( .ip(n5834), .ck(clk), .q(
        \cache_data[7][101] ) );
  dp_1 \cache_data_reg[8][5]  ( .ip(n5802), .ck(clk), .q(\cache_data[8][5] )
         );
  dp_1 \cache_data_reg[8][37]  ( .ip(n5770), .ck(clk), .q(\cache_data[8][37] )
         );
  dp_1 \cache_data_reg[8][69]  ( .ip(n5738), .ck(clk), .q(\cache_data[8][69] )
         );
  dp_1 \cache_data_reg[8][101]  ( .ip(n5706), .ck(clk), .q(
        \cache_data[8][101] ) );
  dp_1 \cache_data_reg[9][5]  ( .ip(n5674), .ck(clk), .q(\cache_data[9][5] )
         );
  dp_1 \cache_data_reg[9][37]  ( .ip(n5642), .ck(clk), .q(\cache_data[9][37] )
         );
  dp_1 \cache_data_reg[9][69]  ( .ip(n5610), .ck(clk), .q(\cache_data[9][69] )
         );
  dp_1 \cache_data_reg[9][101]  ( .ip(n5578), .ck(clk), .q(
        \cache_data[9][101] ) );
  dp_1 \cache_data_reg[10][5]  ( .ip(n5546), .ck(clk), .q(\cache_data[10][5] )
         );
  dp_1 \cache_data_reg[10][37]  ( .ip(n5514), .ck(clk), .q(
        \cache_data[10][37] ) );
  dp_1 \cache_data_reg[10][69]  ( .ip(n5482), .ck(clk), .q(
        \cache_data[10][69] ) );
  dp_1 \cache_data_reg[10][101]  ( .ip(n5450), .ck(clk), .q(
        \cache_data[10][101] ) );
  dp_1 \cache_data_reg[11][5]  ( .ip(n5418), .ck(clk), .q(\cache_data[11][5] )
         );
  dp_1 \cache_data_reg[11][37]  ( .ip(n5386), .ck(clk), .q(
        \cache_data[11][37] ) );
  dp_1 \cache_data_reg[11][69]  ( .ip(n5354), .ck(clk), .q(
        \cache_data[11][69] ) );
  dp_1 \cache_data_reg[11][101]  ( .ip(n5322), .ck(clk), .q(
        \cache_data[11][101] ) );
  dp_1 \cache_data_reg[12][5]  ( .ip(n5290), .ck(clk), .q(\cache_data[12][5] )
         );
  dp_1 \cache_data_reg[12][37]  ( .ip(n5258), .ck(clk), .q(
        \cache_data[12][37] ) );
  dp_1 \cache_data_reg[12][69]  ( .ip(n5226), .ck(clk), .q(
        \cache_data[12][69] ) );
  dp_1 \cache_data_reg[12][101]  ( .ip(n5194), .ck(clk), .q(
        \cache_data[12][101] ) );
  dp_1 \cache_data_reg[13][5]  ( .ip(n5162), .ck(clk), .q(\cache_data[13][5] )
         );
  dp_1 \cache_data_reg[13][37]  ( .ip(n5130), .ck(clk), .q(
        \cache_data[13][37] ) );
  dp_1 \cache_data_reg[13][69]  ( .ip(n5098), .ck(clk), .q(
        \cache_data[13][69] ) );
  dp_1 \cache_data_reg[13][101]  ( .ip(n5066), .ck(clk), .q(
        \cache_data[13][101] ) );
  dp_1 \cache_data_reg[14][5]  ( .ip(n5034), .ck(clk), .q(\cache_data[14][5] )
         );
  dp_1 \cache_data_reg[14][37]  ( .ip(n5002), .ck(clk), .q(
        \cache_data[14][37] ) );
  dp_1 \cache_data_reg[14][69]  ( .ip(n4970), .ck(clk), .q(
        \cache_data[14][69] ) );
  dp_1 \cache_data_reg[14][101]  ( .ip(n4938), .ck(clk), .q(
        \cache_data[14][101] ) );
  dp_1 \cache_data_reg[15][5]  ( .ip(n4906), .ck(clk), .q(\cache_data[15][5] )
         );
  dp_1 \cache_data_reg[15][37]  ( .ip(n4874), .ck(clk), .q(
        \cache_data[15][37] ) );
  dp_1 \cache_data_reg[15][69]  ( .ip(n4842), .ck(clk), .q(
        \cache_data[15][69] ) );
  dp_1 \cache_data_reg[15][101]  ( .ip(n4810), .ck(clk), .q(
        \cache_data[15][101] ) );
  dp_1 \iCache_data_wr_reg[6]  ( .ip(n6857), .ck(clk), .q(iCache_data_wr[6])
         );
  dp_1 \cache_data_reg[0][6]  ( .ip(n6825), .ck(clk), .q(\cache_data[0][6] )
         );
  dp_1 \cache_data_reg[0][38]  ( .ip(n6793), .ck(clk), .q(\cache_data[0][38] )
         );
  dp_1 \cache_data_reg[0][70]  ( .ip(n6761), .ck(clk), .q(\cache_data[0][70] )
         );
  dp_1 \cache_data_reg[0][102]  ( .ip(n6729), .ck(clk), .q(
        \cache_data[0][102] ) );
  dp_1 \cache_data_reg[1][6]  ( .ip(n6697), .ck(clk), .q(\cache_data[1][6] )
         );
  dp_1 \cache_data_reg[1][38]  ( .ip(n6665), .ck(clk), .q(\cache_data[1][38] )
         );
  dp_1 \cache_data_reg[1][70]  ( .ip(n6633), .ck(clk), .q(\cache_data[1][70] )
         );
  dp_1 \cache_data_reg[1][102]  ( .ip(n6601), .ck(clk), .q(
        \cache_data[1][102] ) );
  dp_1 \cache_data_reg[2][6]  ( .ip(n6569), .ck(clk), .q(\cache_data[2][6] )
         );
  dp_1 \cache_data_reg[2][38]  ( .ip(n6537), .ck(clk), .q(\cache_data[2][38] )
         );
  dp_1 \cache_data_reg[2][70]  ( .ip(n6505), .ck(clk), .q(\cache_data[2][70] )
         );
  dp_1 \cache_data_reg[2][102]  ( .ip(n6473), .ck(clk), .q(
        \cache_data[2][102] ) );
  dp_1 \cache_data_reg[3][6]  ( .ip(n6441), .ck(clk), .q(\cache_data[3][6] )
         );
  dp_1 \cache_data_reg[3][38]  ( .ip(n6409), .ck(clk), .q(\cache_data[3][38] )
         );
  dp_1 \cache_data_reg[3][70]  ( .ip(n6377), .ck(clk), .q(\cache_data[3][70] )
         );
  dp_1 \cache_data_reg[3][102]  ( .ip(n6345), .ck(clk), .q(
        \cache_data[3][102] ) );
  dp_1 \cache_data_reg[4][6]  ( .ip(n6313), .ck(clk), .q(\cache_data[4][6] )
         );
  dp_1 \cache_data_reg[4][38]  ( .ip(n6281), .ck(clk), .q(\cache_data[4][38] )
         );
  dp_1 \cache_data_reg[4][70]  ( .ip(n6249), .ck(clk), .q(\cache_data[4][70] )
         );
  dp_1 \cache_data_reg[4][102]  ( .ip(n6217), .ck(clk), .q(
        \cache_data[4][102] ) );
  dp_1 \cache_data_reg[5][6]  ( .ip(n6185), .ck(clk), .q(\cache_data[5][6] )
         );
  dp_1 \cache_data_reg[5][38]  ( .ip(n6153), .ck(clk), .q(\cache_data[5][38] )
         );
  dp_1 \cache_data_reg[5][70]  ( .ip(n6121), .ck(clk), .q(\cache_data[5][70] )
         );
  dp_1 \cache_data_reg[5][102]  ( .ip(n6089), .ck(clk), .q(
        \cache_data[5][102] ) );
  dp_1 \cache_data_reg[6][6]  ( .ip(n6057), .ck(clk), .q(\cache_data[6][6] )
         );
  dp_1 \cache_data_reg[6][38]  ( .ip(n6025), .ck(clk), .q(\cache_data[6][38] )
         );
  dp_1 \cache_data_reg[6][70]  ( .ip(n5993), .ck(clk), .q(\cache_data[6][70] )
         );
  dp_1 \cache_data_reg[6][102]  ( .ip(n5961), .ck(clk), .q(
        \cache_data[6][102] ) );
  dp_1 \cache_data_reg[7][6]  ( .ip(n5929), .ck(clk), .q(\cache_data[7][6] )
         );
  dp_1 \cache_data_reg[7][38]  ( .ip(n5897), .ck(clk), .q(\cache_data[7][38] )
         );
  dp_1 \cache_data_reg[7][70]  ( .ip(n5865), .ck(clk), .q(\cache_data[7][70] )
         );
  dp_1 \cache_data_reg[7][102]  ( .ip(n5833), .ck(clk), .q(
        \cache_data[7][102] ) );
  dp_1 \cache_data_reg[8][6]  ( .ip(n5801), .ck(clk), .q(\cache_data[8][6] )
         );
  dp_1 \cache_data_reg[8][38]  ( .ip(n5769), .ck(clk), .q(\cache_data[8][38] )
         );
  dp_1 \cache_data_reg[8][70]  ( .ip(n5737), .ck(clk), .q(\cache_data[8][70] )
         );
  dp_1 \cache_data_reg[8][102]  ( .ip(n5705), .ck(clk), .q(
        \cache_data[8][102] ) );
  dp_1 \cache_data_reg[9][6]  ( .ip(n5673), .ck(clk), .q(\cache_data[9][6] )
         );
  dp_1 \cache_data_reg[9][38]  ( .ip(n5641), .ck(clk), .q(\cache_data[9][38] )
         );
  dp_1 \cache_data_reg[9][70]  ( .ip(n5609), .ck(clk), .q(\cache_data[9][70] )
         );
  dp_1 \cache_data_reg[9][102]  ( .ip(n5577), .ck(clk), .q(
        \cache_data[9][102] ) );
  dp_1 \cache_data_reg[10][6]  ( .ip(n5545), .ck(clk), .q(\cache_data[10][6] )
         );
  dp_1 \cache_data_reg[10][38]  ( .ip(n5513), .ck(clk), .q(
        \cache_data[10][38] ) );
  dp_1 \cache_data_reg[10][70]  ( .ip(n5481), .ck(clk), .q(
        \cache_data[10][70] ) );
  dp_1 \cache_data_reg[10][102]  ( .ip(n5449), .ck(clk), .q(
        \cache_data[10][102] ) );
  dp_1 \cache_data_reg[11][6]  ( .ip(n5417), .ck(clk), .q(\cache_data[11][6] )
         );
  dp_1 \cache_data_reg[11][38]  ( .ip(n5385), .ck(clk), .q(
        \cache_data[11][38] ) );
  dp_1 \cache_data_reg[11][70]  ( .ip(n5353), .ck(clk), .q(
        \cache_data[11][70] ) );
  dp_1 \cache_data_reg[11][102]  ( .ip(n5321), .ck(clk), .q(
        \cache_data[11][102] ) );
  dp_1 \cache_data_reg[12][6]  ( .ip(n5289), .ck(clk), .q(\cache_data[12][6] )
         );
  dp_1 \cache_data_reg[12][38]  ( .ip(n5257), .ck(clk), .q(
        \cache_data[12][38] ) );
  dp_1 \cache_data_reg[12][70]  ( .ip(n5225), .ck(clk), .q(
        \cache_data[12][70] ) );
  dp_1 \cache_data_reg[12][102]  ( .ip(n5193), .ck(clk), .q(
        \cache_data[12][102] ) );
  dp_1 \cache_data_reg[13][6]  ( .ip(n5161), .ck(clk), .q(\cache_data[13][6] )
         );
  dp_1 \cache_data_reg[13][38]  ( .ip(n5129), .ck(clk), .q(
        \cache_data[13][38] ) );
  dp_1 \cache_data_reg[13][70]  ( .ip(n5097), .ck(clk), .q(
        \cache_data[13][70] ) );
  dp_1 \cache_data_reg[13][102]  ( .ip(n5065), .ck(clk), .q(
        \cache_data[13][102] ) );
  dp_1 \cache_data_reg[14][6]  ( .ip(n5033), .ck(clk), .q(\cache_data[14][6] )
         );
  dp_1 \cache_data_reg[14][38]  ( .ip(n5001), .ck(clk), .q(
        \cache_data[14][38] ) );
  dp_1 \cache_data_reg[14][70]  ( .ip(n4969), .ck(clk), .q(
        \cache_data[14][70] ) );
  dp_1 \cache_data_reg[14][102]  ( .ip(n4937), .ck(clk), .q(
        \cache_data[14][102] ) );
  dp_1 \cache_data_reg[15][6]  ( .ip(n4905), .ck(clk), .q(\cache_data[15][6] )
         );
  dp_1 \cache_data_reg[15][38]  ( .ip(n4873), .ck(clk), .q(
        \cache_data[15][38] ) );
  dp_1 \cache_data_reg[15][70]  ( .ip(n4841), .ck(clk), .q(
        \cache_data[15][70] ) );
  dp_1 \cache_data_reg[15][102]  ( .ip(n4809), .ck(clk), .q(
        \cache_data[15][102] ) );
  dp_1 \iCache_data_wr_reg[7]  ( .ip(n6856), .ck(clk), .q(iCache_data_wr[7])
         );
  dp_1 \cache_data_reg[0][7]  ( .ip(n6824), .ck(clk), .q(\cache_data[0][7] )
         );
  dp_1 \cache_data_reg[0][39]  ( .ip(n6792), .ck(clk), .q(\cache_data[0][39] )
         );
  dp_1 \cache_data_reg[0][71]  ( .ip(n6760), .ck(clk), .q(\cache_data[0][71] )
         );
  dp_1 \cache_data_reg[0][103]  ( .ip(n6728), .ck(clk), .q(
        \cache_data[0][103] ) );
  dp_1 \cache_data_reg[1][7]  ( .ip(n6696), .ck(clk), .q(\cache_data[1][7] )
         );
  dp_1 \cache_data_reg[1][39]  ( .ip(n6664), .ck(clk), .q(\cache_data[1][39] )
         );
  dp_1 \cache_data_reg[1][71]  ( .ip(n6632), .ck(clk), .q(\cache_data[1][71] )
         );
  dp_1 \cache_data_reg[1][103]  ( .ip(n6600), .ck(clk), .q(
        \cache_data[1][103] ) );
  dp_1 \cache_data_reg[2][7]  ( .ip(n6568), .ck(clk), .q(\cache_data[2][7] )
         );
  dp_1 \cache_data_reg[2][39]  ( .ip(n6536), .ck(clk), .q(\cache_data[2][39] )
         );
  dp_1 \cache_data_reg[2][71]  ( .ip(n6504), .ck(clk), .q(\cache_data[2][71] )
         );
  dp_1 \cache_data_reg[2][103]  ( .ip(n6472), .ck(clk), .q(
        \cache_data[2][103] ) );
  dp_1 \cache_data_reg[3][7]  ( .ip(n6440), .ck(clk), .q(\cache_data[3][7] )
         );
  dp_1 \cache_data_reg[3][39]  ( .ip(n6408), .ck(clk), .q(\cache_data[3][39] )
         );
  dp_1 \cache_data_reg[3][71]  ( .ip(n6376), .ck(clk), .q(\cache_data[3][71] )
         );
  dp_1 \cache_data_reg[3][103]  ( .ip(n6344), .ck(clk), .q(
        \cache_data[3][103] ) );
  dp_1 \cache_data_reg[4][7]  ( .ip(n6312), .ck(clk), .q(\cache_data[4][7] )
         );
  dp_1 \cache_data_reg[4][39]  ( .ip(n6280), .ck(clk), .q(\cache_data[4][39] )
         );
  dp_1 \cache_data_reg[4][71]  ( .ip(n6248), .ck(clk), .q(\cache_data[4][71] )
         );
  dp_1 \cache_data_reg[4][103]  ( .ip(n6216), .ck(clk), .q(
        \cache_data[4][103] ) );
  dp_1 \cache_data_reg[5][7]  ( .ip(n6184), .ck(clk), .q(\cache_data[5][7] )
         );
  dp_1 \cache_data_reg[5][39]  ( .ip(n6152), .ck(clk), .q(\cache_data[5][39] )
         );
  dp_1 \cache_data_reg[5][71]  ( .ip(n6120), .ck(clk), .q(\cache_data[5][71] )
         );
  dp_1 \cache_data_reg[5][103]  ( .ip(n6088), .ck(clk), .q(
        \cache_data[5][103] ) );
  dp_1 \cache_data_reg[6][7]  ( .ip(n6056), .ck(clk), .q(\cache_data[6][7] )
         );
  dp_1 \cache_data_reg[6][39]  ( .ip(n6024), .ck(clk), .q(\cache_data[6][39] )
         );
  dp_1 \cache_data_reg[6][71]  ( .ip(n5992), .ck(clk), .q(\cache_data[6][71] )
         );
  dp_1 \cache_data_reg[6][103]  ( .ip(n5960), .ck(clk), .q(
        \cache_data[6][103] ) );
  dp_1 \cache_data_reg[7][7]  ( .ip(n5928), .ck(clk), .q(\cache_data[7][7] )
         );
  dp_1 \cache_data_reg[7][39]  ( .ip(n5896), .ck(clk), .q(\cache_data[7][39] )
         );
  dp_1 \cache_data_reg[7][71]  ( .ip(n5864), .ck(clk), .q(\cache_data[7][71] )
         );
  dp_1 \cache_data_reg[7][103]  ( .ip(n5832), .ck(clk), .q(
        \cache_data[7][103] ) );
  dp_1 \cache_data_reg[8][7]  ( .ip(n5800), .ck(clk), .q(\cache_data[8][7] )
         );
  dp_1 \cache_data_reg[8][39]  ( .ip(n5768), .ck(clk), .q(\cache_data[8][39] )
         );
  dp_1 \cache_data_reg[8][71]  ( .ip(n5736), .ck(clk), .q(\cache_data[8][71] )
         );
  dp_1 \cache_data_reg[8][103]  ( .ip(n5704), .ck(clk), .q(
        \cache_data[8][103] ) );
  dp_1 \cache_data_reg[9][7]  ( .ip(n5672), .ck(clk), .q(\cache_data[9][7] )
         );
  dp_1 \cache_data_reg[9][39]  ( .ip(n5640), .ck(clk), .q(\cache_data[9][39] )
         );
  dp_1 \cache_data_reg[9][71]  ( .ip(n5608), .ck(clk), .q(\cache_data[9][71] )
         );
  dp_1 \cache_data_reg[9][103]  ( .ip(n5576), .ck(clk), .q(
        \cache_data[9][103] ) );
  dp_1 \cache_data_reg[10][7]  ( .ip(n5544), .ck(clk), .q(\cache_data[10][7] )
         );
  dp_1 \cache_data_reg[10][39]  ( .ip(n5512), .ck(clk), .q(
        \cache_data[10][39] ) );
  dp_1 \cache_data_reg[10][71]  ( .ip(n5480), .ck(clk), .q(
        \cache_data[10][71] ) );
  dp_1 \cache_data_reg[10][103]  ( .ip(n5448), .ck(clk), .q(
        \cache_data[10][103] ) );
  dp_1 \cache_data_reg[11][7]  ( .ip(n5416), .ck(clk), .q(\cache_data[11][7] )
         );
  dp_1 \cache_data_reg[11][39]  ( .ip(n5384), .ck(clk), .q(
        \cache_data[11][39] ) );
  dp_1 \cache_data_reg[11][71]  ( .ip(n5352), .ck(clk), .q(
        \cache_data[11][71] ) );
  dp_1 \cache_data_reg[11][103]  ( .ip(n5320), .ck(clk), .q(
        \cache_data[11][103] ) );
  dp_1 \cache_data_reg[12][7]  ( .ip(n5288), .ck(clk), .q(\cache_data[12][7] )
         );
  dp_1 \cache_data_reg[12][39]  ( .ip(n5256), .ck(clk), .q(
        \cache_data[12][39] ) );
  dp_1 \cache_data_reg[12][71]  ( .ip(n5224), .ck(clk), .q(
        \cache_data[12][71] ) );
  dp_1 \cache_data_reg[12][103]  ( .ip(n5192), .ck(clk), .q(
        \cache_data[12][103] ) );
  dp_1 \cache_data_reg[13][7]  ( .ip(n5160), .ck(clk), .q(\cache_data[13][7] )
         );
  dp_1 \cache_data_reg[13][39]  ( .ip(n5128), .ck(clk), .q(
        \cache_data[13][39] ) );
  dp_1 \cache_data_reg[13][71]  ( .ip(n5096), .ck(clk), .q(
        \cache_data[13][71] ) );
  dp_1 \cache_data_reg[13][103]  ( .ip(n5064), .ck(clk), .q(
        \cache_data[13][103] ) );
  dp_1 \cache_data_reg[14][7]  ( .ip(n5032), .ck(clk), .q(\cache_data[14][7] )
         );
  dp_1 \cache_data_reg[14][39]  ( .ip(n5000), .ck(clk), .q(
        \cache_data[14][39] ) );
  dp_1 \cache_data_reg[14][71]  ( .ip(n4968), .ck(clk), .q(
        \cache_data[14][71] ) );
  dp_1 \cache_data_reg[14][103]  ( .ip(n4936), .ck(clk), .q(
        \cache_data[14][103] ) );
  dp_1 \cache_data_reg[15][7]  ( .ip(n4904), .ck(clk), .q(\cache_data[15][7] )
         );
  dp_1 \cache_data_reg[15][39]  ( .ip(n4872), .ck(clk), .q(
        \cache_data[15][39] ) );
  dp_1 \cache_data_reg[15][71]  ( .ip(n4840), .ck(clk), .q(
        \cache_data[15][71] ) );
  dp_1 \cache_data_reg[15][103]  ( .ip(n4808), .ck(clk), .q(
        \cache_data[15][103] ) );
  dp_1 \iCache_data_wr_reg[8]  ( .ip(n6855), .ck(clk), .q(iCache_data_wr[8])
         );
  dp_1 \cache_data_reg[0][8]  ( .ip(n6823), .ck(clk), .q(\cache_data[0][8] )
         );
  dp_1 \cache_data_reg[0][40]  ( .ip(n6791), .ck(clk), .q(\cache_data[0][40] )
         );
  dp_1 \cache_data_reg[0][72]  ( .ip(n6759), .ck(clk), .q(\cache_data[0][72] )
         );
  dp_1 \cache_data_reg[0][104]  ( .ip(n6727), .ck(clk), .q(
        \cache_data[0][104] ) );
  dp_1 \cache_data_reg[1][8]  ( .ip(n6695), .ck(clk), .q(\cache_data[1][8] )
         );
  dp_1 \cache_data_reg[1][40]  ( .ip(n6663), .ck(clk), .q(\cache_data[1][40] )
         );
  dp_1 \cache_data_reg[1][72]  ( .ip(n6631), .ck(clk), .q(\cache_data[1][72] )
         );
  dp_1 \cache_data_reg[1][104]  ( .ip(n6599), .ck(clk), .q(
        \cache_data[1][104] ) );
  dp_1 \cache_data_reg[2][8]  ( .ip(n6567), .ck(clk), .q(\cache_data[2][8] )
         );
  dp_1 \cache_data_reg[2][40]  ( .ip(n6535), .ck(clk), .q(\cache_data[2][40] )
         );
  dp_1 \cache_data_reg[2][72]  ( .ip(n6503), .ck(clk), .q(\cache_data[2][72] )
         );
  dp_1 \cache_data_reg[2][104]  ( .ip(n6471), .ck(clk), .q(
        \cache_data[2][104] ) );
  dp_1 \cache_data_reg[3][8]  ( .ip(n6439), .ck(clk), .q(\cache_data[3][8] )
         );
  dp_1 \cache_data_reg[3][40]  ( .ip(n6407), .ck(clk), .q(\cache_data[3][40] )
         );
  dp_1 \cache_data_reg[3][72]  ( .ip(n6375), .ck(clk), .q(\cache_data[3][72] )
         );
  dp_1 \cache_data_reg[3][104]  ( .ip(n6343), .ck(clk), .q(
        \cache_data[3][104] ) );
  dp_1 \cache_data_reg[4][8]  ( .ip(n6311), .ck(clk), .q(\cache_data[4][8] )
         );
  dp_1 \cache_data_reg[4][40]  ( .ip(n6279), .ck(clk), .q(\cache_data[4][40] )
         );
  dp_1 \cache_data_reg[4][72]  ( .ip(n6247), .ck(clk), .q(\cache_data[4][72] )
         );
  dp_1 \cache_data_reg[4][104]  ( .ip(n6215), .ck(clk), .q(
        \cache_data[4][104] ) );
  dp_1 \cache_data_reg[5][8]  ( .ip(n6183), .ck(clk), .q(\cache_data[5][8] )
         );
  dp_1 \cache_data_reg[5][40]  ( .ip(n6151), .ck(clk), .q(\cache_data[5][40] )
         );
  dp_1 \cache_data_reg[5][72]  ( .ip(n6119), .ck(clk), .q(\cache_data[5][72] )
         );
  dp_1 \cache_data_reg[5][104]  ( .ip(n6087), .ck(clk), .q(
        \cache_data[5][104] ) );
  dp_1 \cache_data_reg[6][8]  ( .ip(n6055), .ck(clk), .q(\cache_data[6][8] )
         );
  dp_1 \cache_data_reg[6][40]  ( .ip(n6023), .ck(clk), .q(\cache_data[6][40] )
         );
  dp_1 \cache_data_reg[6][72]  ( .ip(n5991), .ck(clk), .q(\cache_data[6][72] )
         );
  dp_1 \cache_data_reg[6][104]  ( .ip(n5959), .ck(clk), .q(
        \cache_data[6][104] ) );
  dp_1 \cache_data_reg[7][8]  ( .ip(n5927), .ck(clk), .q(\cache_data[7][8] )
         );
  dp_1 \cache_data_reg[7][40]  ( .ip(n5895), .ck(clk), .q(\cache_data[7][40] )
         );
  dp_1 \cache_data_reg[7][72]  ( .ip(n5863), .ck(clk), .q(\cache_data[7][72] )
         );
  dp_1 \cache_data_reg[7][104]  ( .ip(n5831), .ck(clk), .q(
        \cache_data[7][104] ) );
  dp_1 \cache_data_reg[8][8]  ( .ip(n5799), .ck(clk), .q(\cache_data[8][8] )
         );
  dp_1 \cache_data_reg[8][40]  ( .ip(n5767), .ck(clk), .q(\cache_data[8][40] )
         );
  dp_1 \cache_data_reg[8][72]  ( .ip(n5735), .ck(clk), .q(\cache_data[8][72] )
         );
  dp_1 \cache_data_reg[8][104]  ( .ip(n5703), .ck(clk), .q(
        \cache_data[8][104] ) );
  dp_1 \cache_data_reg[9][8]  ( .ip(n5671), .ck(clk), .q(\cache_data[9][8] )
         );
  dp_1 \cache_data_reg[9][40]  ( .ip(n5639), .ck(clk), .q(\cache_data[9][40] )
         );
  dp_1 \cache_data_reg[9][72]  ( .ip(n5607), .ck(clk), .q(\cache_data[9][72] )
         );
  dp_1 \cache_data_reg[9][104]  ( .ip(n5575), .ck(clk), .q(
        \cache_data[9][104] ) );
  dp_1 \cache_data_reg[10][8]  ( .ip(n5543), .ck(clk), .q(\cache_data[10][8] )
         );
  dp_1 \cache_data_reg[10][40]  ( .ip(n5511), .ck(clk), .q(
        \cache_data[10][40] ) );
  dp_1 \cache_data_reg[10][72]  ( .ip(n5479), .ck(clk), .q(
        \cache_data[10][72] ) );
  dp_1 \cache_data_reg[10][104]  ( .ip(n5447), .ck(clk), .q(
        \cache_data[10][104] ) );
  dp_1 \cache_data_reg[11][8]  ( .ip(n5415), .ck(clk), .q(\cache_data[11][8] )
         );
  dp_1 \cache_data_reg[11][40]  ( .ip(n5383), .ck(clk), .q(
        \cache_data[11][40] ) );
  dp_1 \cache_data_reg[11][72]  ( .ip(n5351), .ck(clk), .q(
        \cache_data[11][72] ) );
  dp_1 \cache_data_reg[11][104]  ( .ip(n5319), .ck(clk), .q(
        \cache_data[11][104] ) );
  dp_1 \cache_data_reg[12][8]  ( .ip(n5287), .ck(clk), .q(\cache_data[12][8] )
         );
  dp_1 \cache_data_reg[12][40]  ( .ip(n5255), .ck(clk), .q(
        \cache_data[12][40] ) );
  dp_1 \cache_data_reg[12][72]  ( .ip(n5223), .ck(clk), .q(
        \cache_data[12][72] ) );
  dp_1 \cache_data_reg[12][104]  ( .ip(n5191), .ck(clk), .q(
        \cache_data[12][104] ) );
  dp_1 \cache_data_reg[13][8]  ( .ip(n5159), .ck(clk), .q(\cache_data[13][8] )
         );
  dp_1 \cache_data_reg[13][40]  ( .ip(n5127), .ck(clk), .q(
        \cache_data[13][40] ) );
  dp_1 \cache_data_reg[13][72]  ( .ip(n5095), .ck(clk), .q(
        \cache_data[13][72] ) );
  dp_1 \cache_data_reg[13][104]  ( .ip(n5063), .ck(clk), .q(
        \cache_data[13][104] ) );
  dp_1 \cache_data_reg[14][8]  ( .ip(n5031), .ck(clk), .q(\cache_data[14][8] )
         );
  dp_1 \cache_data_reg[14][40]  ( .ip(n4999), .ck(clk), .q(
        \cache_data[14][40] ) );
  dp_1 \cache_data_reg[14][72]  ( .ip(n4967), .ck(clk), .q(
        \cache_data[14][72] ) );
  dp_1 \cache_data_reg[14][104]  ( .ip(n4935), .ck(clk), .q(
        \cache_data[14][104] ) );
  dp_1 \cache_data_reg[15][8]  ( .ip(n4903), .ck(clk), .q(\cache_data[15][8] )
         );
  dp_1 \cache_data_reg[15][40]  ( .ip(n4871), .ck(clk), .q(
        \cache_data[15][40] ) );
  dp_1 \cache_data_reg[15][72]  ( .ip(n4839), .ck(clk), .q(
        \cache_data[15][72] ) );
  dp_1 \cache_data_reg[15][104]  ( .ip(n4807), .ck(clk), .q(
        \cache_data[15][104] ) );
  dp_1 \iCache_data_wr_reg[9]  ( .ip(n6854), .ck(clk), .q(iCache_data_wr[9])
         );
  dp_1 \cache_data_reg[0][9]  ( .ip(n6822), .ck(clk), .q(\cache_data[0][9] )
         );
  dp_1 \cache_data_reg[0][41]  ( .ip(n6790), .ck(clk), .q(\cache_data[0][41] )
         );
  dp_1 \cache_data_reg[0][73]  ( .ip(n6758), .ck(clk), .q(\cache_data[0][73] )
         );
  dp_1 \cache_data_reg[0][105]  ( .ip(n6726), .ck(clk), .q(
        \cache_data[0][105] ) );
  dp_1 \cache_data_reg[1][9]  ( .ip(n6694), .ck(clk), .q(\cache_data[1][9] )
         );
  dp_1 \cache_data_reg[1][41]  ( .ip(n6662), .ck(clk), .q(\cache_data[1][41] )
         );
  dp_1 \cache_data_reg[1][73]  ( .ip(n6630), .ck(clk), .q(\cache_data[1][73] )
         );
  dp_1 \cache_data_reg[1][105]  ( .ip(n6598), .ck(clk), .q(
        \cache_data[1][105] ) );
  dp_1 \cache_data_reg[2][9]  ( .ip(n6566), .ck(clk), .q(\cache_data[2][9] )
         );
  dp_1 \cache_data_reg[2][41]  ( .ip(n6534), .ck(clk), .q(\cache_data[2][41] )
         );
  dp_1 \cache_data_reg[2][73]  ( .ip(n6502), .ck(clk), .q(\cache_data[2][73] )
         );
  dp_1 \cache_data_reg[2][105]  ( .ip(n6470), .ck(clk), .q(
        \cache_data[2][105] ) );
  dp_1 \cache_data_reg[3][9]  ( .ip(n6438), .ck(clk), .q(\cache_data[3][9] )
         );
  dp_1 \cache_data_reg[3][41]  ( .ip(n6406), .ck(clk), .q(\cache_data[3][41] )
         );
  dp_1 \cache_data_reg[3][73]  ( .ip(n6374), .ck(clk), .q(\cache_data[3][73] )
         );
  dp_1 \cache_data_reg[3][105]  ( .ip(n6342), .ck(clk), .q(
        \cache_data[3][105] ) );
  dp_1 \cache_data_reg[4][9]  ( .ip(n6310), .ck(clk), .q(\cache_data[4][9] )
         );
  dp_1 \cache_data_reg[4][41]  ( .ip(n6278), .ck(clk), .q(\cache_data[4][41] )
         );
  dp_1 \cache_data_reg[4][73]  ( .ip(n6246), .ck(clk), .q(\cache_data[4][73] )
         );
  dp_1 \cache_data_reg[4][105]  ( .ip(n6214), .ck(clk), .q(
        \cache_data[4][105] ) );
  dp_1 \cache_data_reg[5][9]  ( .ip(n6182), .ck(clk), .q(\cache_data[5][9] )
         );
  dp_1 \cache_data_reg[5][41]  ( .ip(n6150), .ck(clk), .q(\cache_data[5][41] )
         );
  dp_1 \cache_data_reg[5][73]  ( .ip(n6118), .ck(clk), .q(\cache_data[5][73] )
         );
  dp_1 \cache_data_reg[5][105]  ( .ip(n6086), .ck(clk), .q(
        \cache_data[5][105] ) );
  dp_1 \cache_data_reg[6][9]  ( .ip(n6054), .ck(clk), .q(\cache_data[6][9] )
         );
  dp_1 \cache_data_reg[6][41]  ( .ip(n6022), .ck(clk), .q(\cache_data[6][41] )
         );
  dp_1 \cache_data_reg[6][73]  ( .ip(n5990), .ck(clk), .q(\cache_data[6][73] )
         );
  dp_1 \cache_data_reg[6][105]  ( .ip(n5958), .ck(clk), .q(
        \cache_data[6][105] ) );
  dp_1 \cache_data_reg[7][9]  ( .ip(n5926), .ck(clk), .q(\cache_data[7][9] )
         );
  dp_1 \cache_data_reg[7][41]  ( .ip(n5894), .ck(clk), .q(\cache_data[7][41] )
         );
  dp_1 \cache_data_reg[7][73]  ( .ip(n5862), .ck(clk), .q(\cache_data[7][73] )
         );
  dp_1 \cache_data_reg[7][105]  ( .ip(n5830), .ck(clk), .q(
        \cache_data[7][105] ) );
  dp_1 \cache_data_reg[8][9]  ( .ip(n5798), .ck(clk), .q(\cache_data[8][9] )
         );
  dp_1 \cache_data_reg[8][41]  ( .ip(n5766), .ck(clk), .q(\cache_data[8][41] )
         );
  dp_1 \cache_data_reg[8][73]  ( .ip(n5734), .ck(clk), .q(\cache_data[8][73] )
         );
  dp_1 \cache_data_reg[8][105]  ( .ip(n5702), .ck(clk), .q(
        \cache_data[8][105] ) );
  dp_1 \cache_data_reg[9][9]  ( .ip(n5670), .ck(clk), .q(\cache_data[9][9] )
         );
  dp_1 \cache_data_reg[9][41]  ( .ip(n5638), .ck(clk), .q(\cache_data[9][41] )
         );
  dp_1 \cache_data_reg[9][73]  ( .ip(n5606), .ck(clk), .q(\cache_data[9][73] )
         );
  dp_1 \cache_data_reg[9][105]  ( .ip(n5574), .ck(clk), .q(
        \cache_data[9][105] ) );
  dp_1 \cache_data_reg[10][9]  ( .ip(n5542), .ck(clk), .q(\cache_data[10][9] )
         );
  dp_1 \cache_data_reg[10][41]  ( .ip(n5510), .ck(clk), .q(
        \cache_data[10][41] ) );
  dp_1 \cache_data_reg[10][73]  ( .ip(n5478), .ck(clk), .q(
        \cache_data[10][73] ) );
  dp_1 \cache_data_reg[10][105]  ( .ip(n5446), .ck(clk), .q(
        \cache_data[10][105] ) );
  dp_1 \cache_data_reg[11][9]  ( .ip(n5414), .ck(clk), .q(\cache_data[11][9] )
         );
  dp_1 \cache_data_reg[11][41]  ( .ip(n5382), .ck(clk), .q(
        \cache_data[11][41] ) );
  dp_1 \cache_data_reg[11][73]  ( .ip(n5350), .ck(clk), .q(
        \cache_data[11][73] ) );
  dp_1 \cache_data_reg[11][105]  ( .ip(n5318), .ck(clk), .q(
        \cache_data[11][105] ) );
  dp_1 \cache_data_reg[12][9]  ( .ip(n5286), .ck(clk), .q(\cache_data[12][9] )
         );
  dp_1 \cache_data_reg[12][41]  ( .ip(n5254), .ck(clk), .q(
        \cache_data[12][41] ) );
  dp_1 \cache_data_reg[12][73]  ( .ip(n5222), .ck(clk), .q(
        \cache_data[12][73] ) );
  dp_1 \cache_data_reg[12][105]  ( .ip(n5190), .ck(clk), .q(
        \cache_data[12][105] ) );
  dp_1 \cache_data_reg[13][9]  ( .ip(n5158), .ck(clk), .q(\cache_data[13][9] )
         );
  dp_1 \cache_data_reg[13][41]  ( .ip(n5126), .ck(clk), .q(
        \cache_data[13][41] ) );
  dp_1 \cache_data_reg[13][73]  ( .ip(n5094), .ck(clk), .q(
        \cache_data[13][73] ) );
  dp_1 \cache_data_reg[13][105]  ( .ip(n5062), .ck(clk), .q(
        \cache_data[13][105] ) );
  dp_1 \cache_data_reg[14][9]  ( .ip(n5030), .ck(clk), .q(\cache_data[14][9] )
         );
  dp_1 \cache_data_reg[14][41]  ( .ip(n4998), .ck(clk), .q(
        \cache_data[14][41] ) );
  dp_1 \cache_data_reg[14][73]  ( .ip(n4966), .ck(clk), .q(
        \cache_data[14][73] ) );
  dp_1 \cache_data_reg[14][105]  ( .ip(n4934), .ck(clk), .q(
        \cache_data[14][105] ) );
  dp_1 \cache_data_reg[15][9]  ( .ip(n4902), .ck(clk), .q(\cache_data[15][9] )
         );
  dp_1 \cache_data_reg[15][41]  ( .ip(n4870), .ck(clk), .q(
        \cache_data[15][41] ) );
  dp_1 \cache_data_reg[15][73]  ( .ip(n4838), .ck(clk), .q(
        \cache_data[15][73] ) );
  dp_1 \cache_data_reg[15][105]  ( .ip(n4806), .ck(clk), .q(
        \cache_data[15][105] ) );
  dp_1 \iCache_data_wr_reg[10]  ( .ip(n6853), .ck(clk), .q(iCache_data_wr[10])
         );
  dp_1 \cache_data_reg[0][10]  ( .ip(n6821), .ck(clk), .q(\cache_data[0][10] )
         );
  dp_1 \cache_data_reg[0][42]  ( .ip(n6789), .ck(clk), .q(\cache_data[0][42] )
         );
  dp_1 \cache_data_reg[0][74]  ( .ip(n6757), .ck(clk), .q(\cache_data[0][74] )
         );
  dp_1 \cache_data_reg[0][106]  ( .ip(n6725), .ck(clk), .q(
        \cache_data[0][106] ) );
  dp_1 \cache_data_reg[1][10]  ( .ip(n6693), .ck(clk), .q(\cache_data[1][10] )
         );
  dp_1 \cache_data_reg[1][42]  ( .ip(n6661), .ck(clk), .q(\cache_data[1][42] )
         );
  dp_1 \cache_data_reg[1][74]  ( .ip(n6629), .ck(clk), .q(\cache_data[1][74] )
         );
  dp_1 \cache_data_reg[1][106]  ( .ip(n6597), .ck(clk), .q(
        \cache_data[1][106] ) );
  dp_1 \cache_data_reg[2][10]  ( .ip(n6565), .ck(clk), .q(\cache_data[2][10] )
         );
  dp_1 \cache_data_reg[2][42]  ( .ip(n6533), .ck(clk), .q(\cache_data[2][42] )
         );
  dp_1 \cache_data_reg[2][74]  ( .ip(n6501), .ck(clk), .q(\cache_data[2][74] )
         );
  dp_1 \cache_data_reg[2][106]  ( .ip(n6469), .ck(clk), .q(
        \cache_data[2][106] ) );
  dp_1 \cache_data_reg[3][10]  ( .ip(n6437), .ck(clk), .q(\cache_data[3][10] )
         );
  dp_1 \cache_data_reg[3][42]  ( .ip(n6405), .ck(clk), .q(\cache_data[3][42] )
         );
  dp_1 \cache_data_reg[3][74]  ( .ip(n6373), .ck(clk), .q(\cache_data[3][74] )
         );
  dp_1 \cache_data_reg[3][106]  ( .ip(n6341), .ck(clk), .q(
        \cache_data[3][106] ) );
  dp_1 \cache_data_reg[4][10]  ( .ip(n6309), .ck(clk), .q(\cache_data[4][10] )
         );
  dp_1 \cache_data_reg[4][42]  ( .ip(n6277), .ck(clk), .q(\cache_data[4][42] )
         );
  dp_1 \cache_data_reg[4][74]  ( .ip(n6245), .ck(clk), .q(\cache_data[4][74] )
         );
  dp_1 \cache_data_reg[4][106]  ( .ip(n6213), .ck(clk), .q(
        \cache_data[4][106] ) );
  dp_1 \cache_data_reg[5][10]  ( .ip(n6181), .ck(clk), .q(\cache_data[5][10] )
         );
  dp_1 \cache_data_reg[5][42]  ( .ip(n6149), .ck(clk), .q(\cache_data[5][42] )
         );
  dp_1 \cache_data_reg[5][74]  ( .ip(n6117), .ck(clk), .q(\cache_data[5][74] )
         );
  dp_1 \cache_data_reg[5][106]  ( .ip(n6085), .ck(clk), .q(
        \cache_data[5][106] ) );
  dp_1 \cache_data_reg[6][10]  ( .ip(n6053), .ck(clk), .q(\cache_data[6][10] )
         );
  dp_1 \cache_data_reg[6][42]  ( .ip(n6021), .ck(clk), .q(\cache_data[6][42] )
         );
  dp_1 \cache_data_reg[6][74]  ( .ip(n5989), .ck(clk), .q(\cache_data[6][74] )
         );
  dp_1 \cache_data_reg[6][106]  ( .ip(n5957), .ck(clk), .q(
        \cache_data[6][106] ) );
  dp_1 \cache_data_reg[7][10]  ( .ip(n5925), .ck(clk), .q(\cache_data[7][10] )
         );
  dp_1 \cache_data_reg[7][42]  ( .ip(n5893), .ck(clk), .q(\cache_data[7][42] )
         );
  dp_1 \cache_data_reg[7][74]  ( .ip(n5861), .ck(clk), .q(\cache_data[7][74] )
         );
  dp_1 \cache_data_reg[7][106]  ( .ip(n5829), .ck(clk), .q(
        \cache_data[7][106] ) );
  dp_1 \cache_data_reg[8][10]  ( .ip(n5797), .ck(clk), .q(\cache_data[8][10] )
         );
  dp_1 \cache_data_reg[8][42]  ( .ip(n5765), .ck(clk), .q(\cache_data[8][42] )
         );
  dp_1 \cache_data_reg[8][74]  ( .ip(n5733), .ck(clk), .q(\cache_data[8][74] )
         );
  dp_1 \cache_data_reg[8][106]  ( .ip(n5701), .ck(clk), .q(
        \cache_data[8][106] ) );
  dp_1 \cache_data_reg[9][10]  ( .ip(n5669), .ck(clk), .q(\cache_data[9][10] )
         );
  dp_1 \cache_data_reg[9][42]  ( .ip(n5637), .ck(clk), .q(\cache_data[9][42] )
         );
  dp_1 \cache_data_reg[9][74]  ( .ip(n5605), .ck(clk), .q(\cache_data[9][74] )
         );
  dp_1 \cache_data_reg[9][106]  ( .ip(n5573), .ck(clk), .q(
        \cache_data[9][106] ) );
  dp_1 \cache_data_reg[10][10]  ( .ip(n5541), .ck(clk), .q(
        \cache_data[10][10] ) );
  dp_1 \cache_data_reg[10][42]  ( .ip(n5509), .ck(clk), .q(
        \cache_data[10][42] ) );
  dp_1 \cache_data_reg[10][74]  ( .ip(n5477), .ck(clk), .q(
        \cache_data[10][74] ) );
  dp_1 \cache_data_reg[10][106]  ( .ip(n5445), .ck(clk), .q(
        \cache_data[10][106] ) );
  dp_1 \cache_data_reg[11][10]  ( .ip(n5413), .ck(clk), .q(
        \cache_data[11][10] ) );
  dp_1 \cache_data_reg[11][42]  ( .ip(n5381), .ck(clk), .q(
        \cache_data[11][42] ) );
  dp_1 \cache_data_reg[11][74]  ( .ip(n5349), .ck(clk), .q(
        \cache_data[11][74] ) );
  dp_1 \cache_data_reg[11][106]  ( .ip(n5317), .ck(clk), .q(
        \cache_data[11][106] ) );
  dp_1 \cache_data_reg[12][10]  ( .ip(n5285), .ck(clk), .q(
        \cache_data[12][10] ) );
  dp_1 \cache_data_reg[12][42]  ( .ip(n5253), .ck(clk), .q(
        \cache_data[12][42] ) );
  dp_1 \cache_data_reg[12][74]  ( .ip(n5221), .ck(clk), .q(
        \cache_data[12][74] ) );
  dp_1 \cache_data_reg[12][106]  ( .ip(n5189), .ck(clk), .q(
        \cache_data[12][106] ) );
  dp_1 \cache_data_reg[13][10]  ( .ip(n5157), .ck(clk), .q(
        \cache_data[13][10] ) );
  dp_1 \cache_data_reg[13][42]  ( .ip(n5125), .ck(clk), .q(
        \cache_data[13][42] ) );
  dp_1 \cache_data_reg[13][74]  ( .ip(n5093), .ck(clk), .q(
        \cache_data[13][74] ) );
  dp_1 \cache_data_reg[13][106]  ( .ip(n5061), .ck(clk), .q(
        \cache_data[13][106] ) );
  dp_1 \cache_data_reg[14][10]  ( .ip(n5029), .ck(clk), .q(
        \cache_data[14][10] ) );
  dp_1 \cache_data_reg[14][42]  ( .ip(n4997), .ck(clk), .q(
        \cache_data[14][42] ) );
  dp_1 \cache_data_reg[14][74]  ( .ip(n4965), .ck(clk), .q(
        \cache_data[14][74] ) );
  dp_1 \cache_data_reg[14][106]  ( .ip(n4933), .ck(clk), .q(
        \cache_data[14][106] ) );
  dp_1 \cache_data_reg[15][10]  ( .ip(n4901), .ck(clk), .q(
        \cache_data[15][10] ) );
  dp_1 \cache_data_reg[15][42]  ( .ip(n4869), .ck(clk), .q(
        \cache_data[15][42] ) );
  dp_1 \cache_data_reg[15][74]  ( .ip(n4837), .ck(clk), .q(
        \cache_data[15][74] ) );
  dp_1 \cache_data_reg[15][106]  ( .ip(n4805), .ck(clk), .q(
        \cache_data[15][106] ) );
  dp_1 \iCache_data_wr_reg[11]  ( .ip(n6852), .ck(clk), .q(iCache_data_wr[11])
         );
  dp_1 \cache_data_reg[0][11]  ( .ip(n6820), .ck(clk), .q(\cache_data[0][11] )
         );
  dp_1 \cache_data_reg[0][43]  ( .ip(n6788), .ck(clk), .q(\cache_data[0][43] )
         );
  dp_1 \cache_data_reg[0][75]  ( .ip(n6756), .ck(clk), .q(\cache_data[0][75] )
         );
  dp_1 \cache_data_reg[0][107]  ( .ip(n6724), .ck(clk), .q(
        \cache_data[0][107] ) );
  dp_1 \cache_data_reg[1][11]  ( .ip(n6692), .ck(clk), .q(\cache_data[1][11] )
         );
  dp_1 \cache_data_reg[1][43]  ( .ip(n6660), .ck(clk), .q(\cache_data[1][43] )
         );
  dp_1 \cache_data_reg[1][75]  ( .ip(n6628), .ck(clk), .q(\cache_data[1][75] )
         );
  dp_1 \cache_data_reg[1][107]  ( .ip(n6596), .ck(clk), .q(
        \cache_data[1][107] ) );
  dp_1 \cache_data_reg[2][11]  ( .ip(n6564), .ck(clk), .q(\cache_data[2][11] )
         );
  dp_1 \cache_data_reg[2][43]  ( .ip(n6532), .ck(clk), .q(\cache_data[2][43] )
         );
  dp_1 \cache_data_reg[2][75]  ( .ip(n6500), .ck(clk), .q(\cache_data[2][75] )
         );
  dp_1 \cache_data_reg[2][107]  ( .ip(n6468), .ck(clk), .q(
        \cache_data[2][107] ) );
  dp_1 \cache_data_reg[3][11]  ( .ip(n6436), .ck(clk), .q(\cache_data[3][11] )
         );
  dp_1 \cache_data_reg[3][43]  ( .ip(n6404), .ck(clk), .q(\cache_data[3][43] )
         );
  dp_1 \cache_data_reg[3][75]  ( .ip(n6372), .ck(clk), .q(\cache_data[3][75] )
         );
  dp_1 \cache_data_reg[3][107]  ( .ip(n6340), .ck(clk), .q(
        \cache_data[3][107] ) );
  dp_1 \cache_data_reg[4][11]  ( .ip(n6308), .ck(clk), .q(\cache_data[4][11] )
         );
  dp_1 \cache_data_reg[4][43]  ( .ip(n6276), .ck(clk), .q(\cache_data[4][43] )
         );
  dp_1 \cache_data_reg[4][75]  ( .ip(n6244), .ck(clk), .q(\cache_data[4][75] )
         );
  dp_1 \cache_data_reg[4][107]  ( .ip(n6212), .ck(clk), .q(
        \cache_data[4][107] ) );
  dp_1 \cache_data_reg[5][11]  ( .ip(n6180), .ck(clk), .q(\cache_data[5][11] )
         );
  dp_1 \cache_data_reg[5][43]  ( .ip(n6148), .ck(clk), .q(\cache_data[5][43] )
         );
  dp_1 \cache_data_reg[5][75]  ( .ip(n6116), .ck(clk), .q(\cache_data[5][75] )
         );
  dp_1 \cache_data_reg[5][107]  ( .ip(n6084), .ck(clk), .q(
        \cache_data[5][107] ) );
  dp_1 \cache_data_reg[6][11]  ( .ip(n6052), .ck(clk), .q(\cache_data[6][11] )
         );
  dp_1 \cache_data_reg[6][43]  ( .ip(n6020), .ck(clk), .q(\cache_data[6][43] )
         );
  dp_1 \cache_data_reg[6][75]  ( .ip(n5988), .ck(clk), .q(\cache_data[6][75] )
         );
  dp_1 \cache_data_reg[6][107]  ( .ip(n5956), .ck(clk), .q(
        \cache_data[6][107] ) );
  dp_1 \cache_data_reg[7][11]  ( .ip(n5924), .ck(clk), .q(\cache_data[7][11] )
         );
  dp_1 \cache_data_reg[7][43]  ( .ip(n5892), .ck(clk), .q(\cache_data[7][43] )
         );
  dp_1 \cache_data_reg[7][75]  ( .ip(n5860), .ck(clk), .q(\cache_data[7][75] )
         );
  dp_1 \cache_data_reg[7][107]  ( .ip(n5828), .ck(clk), .q(
        \cache_data[7][107] ) );
  dp_1 \cache_data_reg[8][11]  ( .ip(n5796), .ck(clk), .q(\cache_data[8][11] )
         );
  dp_1 \cache_data_reg[8][43]  ( .ip(n5764), .ck(clk), .q(\cache_data[8][43] )
         );
  dp_1 \cache_data_reg[8][75]  ( .ip(n5732), .ck(clk), .q(\cache_data[8][75] )
         );
  dp_1 \cache_data_reg[8][107]  ( .ip(n5700), .ck(clk), .q(
        \cache_data[8][107] ) );
  dp_1 \cache_data_reg[9][11]  ( .ip(n5668), .ck(clk), .q(\cache_data[9][11] )
         );
  dp_1 \cache_data_reg[9][43]  ( .ip(n5636), .ck(clk), .q(\cache_data[9][43] )
         );
  dp_1 \cache_data_reg[9][75]  ( .ip(n5604), .ck(clk), .q(\cache_data[9][75] )
         );
  dp_1 \cache_data_reg[9][107]  ( .ip(n5572), .ck(clk), .q(
        \cache_data[9][107] ) );
  dp_1 \cache_data_reg[10][11]  ( .ip(n5540), .ck(clk), .q(
        \cache_data[10][11] ) );
  dp_1 \cache_data_reg[10][43]  ( .ip(n5508), .ck(clk), .q(
        \cache_data[10][43] ) );
  dp_1 \cache_data_reg[10][75]  ( .ip(n5476), .ck(clk), .q(
        \cache_data[10][75] ) );
  dp_1 \cache_data_reg[10][107]  ( .ip(n5444), .ck(clk), .q(
        \cache_data[10][107] ) );
  dp_1 \cache_data_reg[11][11]  ( .ip(n5412), .ck(clk), .q(
        \cache_data[11][11] ) );
  dp_1 \cache_data_reg[11][43]  ( .ip(n5380), .ck(clk), .q(
        \cache_data[11][43] ) );
  dp_1 \cache_data_reg[11][75]  ( .ip(n5348), .ck(clk), .q(
        \cache_data[11][75] ) );
  dp_1 \cache_data_reg[11][107]  ( .ip(n5316), .ck(clk), .q(
        \cache_data[11][107] ) );
  dp_1 \cache_data_reg[12][11]  ( .ip(n5284), .ck(clk), .q(
        \cache_data[12][11] ) );
  dp_1 \cache_data_reg[12][43]  ( .ip(n5252), .ck(clk), .q(
        \cache_data[12][43] ) );
  dp_1 \cache_data_reg[12][75]  ( .ip(n5220), .ck(clk), .q(
        \cache_data[12][75] ) );
  dp_1 \cache_data_reg[12][107]  ( .ip(n5188), .ck(clk), .q(
        \cache_data[12][107] ) );
  dp_1 \cache_data_reg[13][11]  ( .ip(n5156), .ck(clk), .q(
        \cache_data[13][11] ) );
  dp_1 \cache_data_reg[13][43]  ( .ip(n5124), .ck(clk), .q(
        \cache_data[13][43] ) );
  dp_1 \cache_data_reg[13][75]  ( .ip(n5092), .ck(clk), .q(
        \cache_data[13][75] ) );
  dp_1 \cache_data_reg[13][107]  ( .ip(n5060), .ck(clk), .q(
        \cache_data[13][107] ) );
  dp_1 \cache_data_reg[14][11]  ( .ip(n5028), .ck(clk), .q(
        \cache_data[14][11] ) );
  dp_1 \cache_data_reg[14][43]  ( .ip(n4996), .ck(clk), .q(
        \cache_data[14][43] ) );
  dp_1 \cache_data_reg[14][75]  ( .ip(n4964), .ck(clk), .q(
        \cache_data[14][75] ) );
  dp_1 \cache_data_reg[14][107]  ( .ip(n4932), .ck(clk), .q(
        \cache_data[14][107] ) );
  dp_1 \cache_data_reg[15][11]  ( .ip(n4900), .ck(clk), .q(
        \cache_data[15][11] ) );
  dp_1 \cache_data_reg[15][43]  ( .ip(n4868), .ck(clk), .q(
        \cache_data[15][43] ) );
  dp_1 \cache_data_reg[15][75]  ( .ip(n4836), .ck(clk), .q(
        \cache_data[15][75] ) );
  dp_1 \cache_data_reg[15][107]  ( .ip(n4804), .ck(clk), .q(
        \cache_data[15][107] ) );
  dp_1 \iCache_data_wr_reg[12]  ( .ip(n6851), .ck(clk), .q(iCache_data_wr[12])
         );
  dp_1 \cache_data_reg[0][12]  ( .ip(n6819), .ck(clk), .q(\cache_data[0][12] )
         );
  dp_1 \cache_data_reg[0][44]  ( .ip(n6787), .ck(clk), .q(\cache_data[0][44] )
         );
  dp_1 \cache_data_reg[0][76]  ( .ip(n6755), .ck(clk), .q(\cache_data[0][76] )
         );
  dp_1 \cache_data_reg[0][108]  ( .ip(n6723), .ck(clk), .q(
        \cache_data[0][108] ) );
  dp_1 \cache_data_reg[1][12]  ( .ip(n6691), .ck(clk), .q(\cache_data[1][12] )
         );
  dp_1 \cache_data_reg[1][44]  ( .ip(n6659), .ck(clk), .q(\cache_data[1][44] )
         );
  dp_1 \cache_data_reg[1][76]  ( .ip(n6627), .ck(clk), .q(\cache_data[1][76] )
         );
  dp_1 \cache_data_reg[1][108]  ( .ip(n6595), .ck(clk), .q(
        \cache_data[1][108] ) );
  dp_1 \cache_data_reg[2][12]  ( .ip(n6563), .ck(clk), .q(\cache_data[2][12] )
         );
  dp_1 \cache_data_reg[2][44]  ( .ip(n6531), .ck(clk), .q(\cache_data[2][44] )
         );
  dp_1 \cache_data_reg[2][76]  ( .ip(n6499), .ck(clk), .q(\cache_data[2][76] )
         );
  dp_1 \cache_data_reg[2][108]  ( .ip(n6467), .ck(clk), .q(
        \cache_data[2][108] ) );
  dp_1 \cache_data_reg[3][12]  ( .ip(n6435), .ck(clk), .q(\cache_data[3][12] )
         );
  dp_1 \cache_data_reg[3][44]  ( .ip(n6403), .ck(clk), .q(\cache_data[3][44] )
         );
  dp_1 \cache_data_reg[3][76]  ( .ip(n6371), .ck(clk), .q(\cache_data[3][76] )
         );
  dp_1 \cache_data_reg[3][108]  ( .ip(n6339), .ck(clk), .q(
        \cache_data[3][108] ) );
  dp_1 \cache_data_reg[4][12]  ( .ip(n6307), .ck(clk), .q(\cache_data[4][12] )
         );
  dp_1 \cache_data_reg[4][44]  ( .ip(n6275), .ck(clk), .q(\cache_data[4][44] )
         );
  dp_1 \cache_data_reg[4][76]  ( .ip(n6243), .ck(clk), .q(\cache_data[4][76] )
         );
  dp_1 \cache_data_reg[4][108]  ( .ip(n6211), .ck(clk), .q(
        \cache_data[4][108] ) );
  dp_1 \cache_data_reg[5][12]  ( .ip(n6179), .ck(clk), .q(\cache_data[5][12] )
         );
  dp_1 \cache_data_reg[5][44]  ( .ip(n6147), .ck(clk), .q(\cache_data[5][44] )
         );
  dp_1 \cache_data_reg[5][76]  ( .ip(n6115), .ck(clk), .q(\cache_data[5][76] )
         );
  dp_1 \cache_data_reg[5][108]  ( .ip(n6083), .ck(clk), .q(
        \cache_data[5][108] ) );
  dp_1 \cache_data_reg[6][12]  ( .ip(n6051), .ck(clk), .q(\cache_data[6][12] )
         );
  dp_1 \cache_data_reg[6][44]  ( .ip(n6019), .ck(clk), .q(\cache_data[6][44] )
         );
  dp_1 \cache_data_reg[6][76]  ( .ip(n5987), .ck(clk), .q(\cache_data[6][76] )
         );
  dp_1 \cache_data_reg[6][108]  ( .ip(n5955), .ck(clk), .q(
        \cache_data[6][108] ) );
  dp_1 \cache_data_reg[7][12]  ( .ip(n5923), .ck(clk), .q(\cache_data[7][12] )
         );
  dp_1 \cache_data_reg[7][44]  ( .ip(n5891), .ck(clk), .q(\cache_data[7][44] )
         );
  dp_1 \cache_data_reg[7][76]  ( .ip(n5859), .ck(clk), .q(\cache_data[7][76] )
         );
  dp_1 \cache_data_reg[7][108]  ( .ip(n5827), .ck(clk), .q(
        \cache_data[7][108] ) );
  dp_1 \cache_data_reg[8][12]  ( .ip(n5795), .ck(clk), .q(\cache_data[8][12] )
         );
  dp_1 \cache_data_reg[8][44]  ( .ip(n5763), .ck(clk), .q(\cache_data[8][44] )
         );
  dp_1 \cache_data_reg[8][76]  ( .ip(n5731), .ck(clk), .q(\cache_data[8][76] )
         );
  dp_1 \cache_data_reg[8][108]  ( .ip(n5699), .ck(clk), .q(
        \cache_data[8][108] ) );
  dp_1 \cache_data_reg[9][12]  ( .ip(n5667), .ck(clk), .q(\cache_data[9][12] )
         );
  dp_1 \cache_data_reg[9][44]  ( .ip(n5635), .ck(clk), .q(\cache_data[9][44] )
         );
  dp_1 \cache_data_reg[9][76]  ( .ip(n5603), .ck(clk), .q(\cache_data[9][76] )
         );
  dp_1 \cache_data_reg[9][108]  ( .ip(n5571), .ck(clk), .q(
        \cache_data[9][108] ) );
  dp_1 \cache_data_reg[10][12]  ( .ip(n5539), .ck(clk), .q(
        \cache_data[10][12] ) );
  dp_1 \cache_data_reg[10][44]  ( .ip(n5507), .ck(clk), .q(
        \cache_data[10][44] ) );
  dp_1 \cache_data_reg[10][76]  ( .ip(n5475), .ck(clk), .q(
        \cache_data[10][76] ) );
  dp_1 \cache_data_reg[10][108]  ( .ip(n5443), .ck(clk), .q(
        \cache_data[10][108] ) );
  dp_1 \cache_data_reg[11][12]  ( .ip(n5411), .ck(clk), .q(
        \cache_data[11][12] ) );
  dp_1 \cache_data_reg[11][44]  ( .ip(n5379), .ck(clk), .q(
        \cache_data[11][44] ) );
  dp_1 \cache_data_reg[11][76]  ( .ip(n5347), .ck(clk), .q(
        \cache_data[11][76] ) );
  dp_1 \cache_data_reg[11][108]  ( .ip(n5315), .ck(clk), .q(
        \cache_data[11][108] ) );
  dp_1 \cache_data_reg[12][12]  ( .ip(n5283), .ck(clk), .q(
        \cache_data[12][12] ) );
  dp_1 \cache_data_reg[12][44]  ( .ip(n5251), .ck(clk), .q(
        \cache_data[12][44] ) );
  dp_1 \cache_data_reg[12][76]  ( .ip(n5219), .ck(clk), .q(
        \cache_data[12][76] ) );
  dp_1 \cache_data_reg[12][108]  ( .ip(n5187), .ck(clk), .q(
        \cache_data[12][108] ) );
  dp_1 \cache_data_reg[13][12]  ( .ip(n5155), .ck(clk), .q(
        \cache_data[13][12] ) );
  dp_1 \cache_data_reg[13][44]  ( .ip(n5123), .ck(clk), .q(
        \cache_data[13][44] ) );
  dp_1 \cache_data_reg[13][76]  ( .ip(n5091), .ck(clk), .q(
        \cache_data[13][76] ) );
  dp_1 \cache_data_reg[13][108]  ( .ip(n5059), .ck(clk), .q(
        \cache_data[13][108] ) );
  dp_1 \cache_data_reg[14][12]  ( .ip(n5027), .ck(clk), .q(
        \cache_data[14][12] ) );
  dp_1 \cache_data_reg[14][44]  ( .ip(n4995), .ck(clk), .q(
        \cache_data[14][44] ) );
  dp_1 \cache_data_reg[14][76]  ( .ip(n4963), .ck(clk), .q(
        \cache_data[14][76] ) );
  dp_1 \cache_data_reg[14][108]  ( .ip(n4931), .ck(clk), .q(
        \cache_data[14][108] ) );
  dp_1 \cache_data_reg[15][12]  ( .ip(n4899), .ck(clk), .q(
        \cache_data[15][12] ) );
  dp_1 \cache_data_reg[15][44]  ( .ip(n4867), .ck(clk), .q(
        \cache_data[15][44] ) );
  dp_1 \cache_data_reg[15][76]  ( .ip(n4835), .ck(clk), .q(
        \cache_data[15][76] ) );
  dp_1 \cache_data_reg[15][108]  ( .ip(n4803), .ck(clk), .q(
        \cache_data[15][108] ) );
  dp_1 \iCache_data_wr_reg[13]  ( .ip(n6850), .ck(clk), .q(iCache_data_wr[13])
         );
  dp_1 \cache_data_reg[0][13]  ( .ip(n6818), .ck(clk), .q(\cache_data[0][13] )
         );
  dp_1 \cache_data_reg[0][45]  ( .ip(n6786), .ck(clk), .q(\cache_data[0][45] )
         );
  dp_1 \cache_data_reg[0][77]  ( .ip(n6754), .ck(clk), .q(\cache_data[0][77] )
         );
  dp_1 \cache_data_reg[0][109]  ( .ip(n6722), .ck(clk), .q(
        \cache_data[0][109] ) );
  dp_1 \cache_data_reg[1][13]  ( .ip(n6690), .ck(clk), .q(\cache_data[1][13] )
         );
  dp_1 \cache_data_reg[1][45]  ( .ip(n6658), .ck(clk), .q(\cache_data[1][45] )
         );
  dp_1 \cache_data_reg[1][77]  ( .ip(n6626), .ck(clk), .q(\cache_data[1][77] )
         );
  dp_1 \cache_data_reg[1][109]  ( .ip(n6594), .ck(clk), .q(
        \cache_data[1][109] ) );
  dp_1 \cache_data_reg[2][13]  ( .ip(n6562), .ck(clk), .q(\cache_data[2][13] )
         );
  dp_1 \cache_data_reg[2][45]  ( .ip(n6530), .ck(clk), .q(\cache_data[2][45] )
         );
  dp_1 \cache_data_reg[2][77]  ( .ip(n6498), .ck(clk), .q(\cache_data[2][77] )
         );
  dp_1 \cache_data_reg[2][109]  ( .ip(n6466), .ck(clk), .q(
        \cache_data[2][109] ) );
  dp_1 \cache_data_reg[3][13]  ( .ip(n6434), .ck(clk), .q(\cache_data[3][13] )
         );
  dp_1 \cache_data_reg[3][45]  ( .ip(n6402), .ck(clk), .q(\cache_data[3][45] )
         );
  dp_1 \cache_data_reg[3][77]  ( .ip(n6370), .ck(clk), .q(\cache_data[3][77] )
         );
  dp_1 \cache_data_reg[3][109]  ( .ip(n6338), .ck(clk), .q(
        \cache_data[3][109] ) );
  dp_1 \cache_data_reg[4][13]  ( .ip(n6306), .ck(clk), .q(\cache_data[4][13] )
         );
  dp_1 \cache_data_reg[4][45]  ( .ip(n6274), .ck(clk), .q(\cache_data[4][45] )
         );
  dp_1 \cache_data_reg[4][77]  ( .ip(n6242), .ck(clk), .q(\cache_data[4][77] )
         );
  dp_1 \cache_data_reg[4][109]  ( .ip(n6210), .ck(clk), .q(
        \cache_data[4][109] ) );
  dp_1 \cache_data_reg[5][13]  ( .ip(n6178), .ck(clk), .q(\cache_data[5][13] )
         );
  dp_1 \cache_data_reg[5][45]  ( .ip(n6146), .ck(clk), .q(\cache_data[5][45] )
         );
  dp_1 \cache_data_reg[5][77]  ( .ip(n6114), .ck(clk), .q(\cache_data[5][77] )
         );
  dp_1 \cache_data_reg[5][109]  ( .ip(n6082), .ck(clk), .q(
        \cache_data[5][109] ) );
  dp_1 \cache_data_reg[6][13]  ( .ip(n6050), .ck(clk), .q(\cache_data[6][13] )
         );
  dp_1 \cache_data_reg[6][45]  ( .ip(n6018), .ck(clk), .q(\cache_data[6][45] )
         );
  dp_1 \cache_data_reg[6][77]  ( .ip(n5986), .ck(clk), .q(\cache_data[6][77] )
         );
  dp_1 \cache_data_reg[6][109]  ( .ip(n5954), .ck(clk), .q(
        \cache_data[6][109] ) );
  dp_1 \cache_data_reg[7][13]  ( .ip(n5922), .ck(clk), .q(\cache_data[7][13] )
         );
  dp_1 \cache_data_reg[7][45]  ( .ip(n5890), .ck(clk), .q(\cache_data[7][45] )
         );
  dp_1 \cache_data_reg[7][77]  ( .ip(n5858), .ck(clk), .q(\cache_data[7][77] )
         );
  dp_1 \cache_data_reg[7][109]  ( .ip(n5826), .ck(clk), .q(
        \cache_data[7][109] ) );
  dp_1 \cache_data_reg[8][13]  ( .ip(n5794), .ck(clk), .q(\cache_data[8][13] )
         );
  dp_1 \cache_data_reg[8][45]  ( .ip(n5762), .ck(clk), .q(\cache_data[8][45] )
         );
  dp_1 \cache_data_reg[8][77]  ( .ip(n5730), .ck(clk), .q(\cache_data[8][77] )
         );
  dp_1 \cache_data_reg[8][109]  ( .ip(n5698), .ck(clk), .q(
        \cache_data[8][109] ) );
  dp_1 \cache_data_reg[9][13]  ( .ip(n5666), .ck(clk), .q(\cache_data[9][13] )
         );
  dp_1 \cache_data_reg[9][45]  ( .ip(n5634), .ck(clk), .q(\cache_data[9][45] )
         );
  dp_1 \cache_data_reg[9][77]  ( .ip(n5602), .ck(clk), .q(\cache_data[9][77] )
         );
  dp_1 \cache_data_reg[9][109]  ( .ip(n5570), .ck(clk), .q(
        \cache_data[9][109] ) );
  dp_1 \cache_data_reg[10][13]  ( .ip(n5538), .ck(clk), .q(
        \cache_data[10][13] ) );
  dp_1 \cache_data_reg[10][45]  ( .ip(n5506), .ck(clk), .q(
        \cache_data[10][45] ) );
  dp_1 \cache_data_reg[10][77]  ( .ip(n5474), .ck(clk), .q(
        \cache_data[10][77] ) );
  dp_1 \cache_data_reg[10][109]  ( .ip(n5442), .ck(clk), .q(
        \cache_data[10][109] ) );
  dp_1 \cache_data_reg[11][13]  ( .ip(n5410), .ck(clk), .q(
        \cache_data[11][13] ) );
  dp_1 \cache_data_reg[11][45]  ( .ip(n5378), .ck(clk), .q(
        \cache_data[11][45] ) );
  dp_1 \cache_data_reg[11][77]  ( .ip(n5346), .ck(clk), .q(
        \cache_data[11][77] ) );
  dp_1 \cache_data_reg[11][109]  ( .ip(n5314), .ck(clk), .q(
        \cache_data[11][109] ) );
  dp_1 \cache_data_reg[12][13]  ( .ip(n5282), .ck(clk), .q(
        \cache_data[12][13] ) );
  dp_1 \cache_data_reg[12][45]  ( .ip(n5250), .ck(clk), .q(
        \cache_data[12][45] ) );
  dp_1 \cache_data_reg[12][77]  ( .ip(n5218), .ck(clk), .q(
        \cache_data[12][77] ) );
  dp_1 \cache_data_reg[12][109]  ( .ip(n5186), .ck(clk), .q(
        \cache_data[12][109] ) );
  dp_1 \cache_data_reg[13][13]  ( .ip(n5154), .ck(clk), .q(
        \cache_data[13][13] ) );
  dp_1 \cache_data_reg[13][45]  ( .ip(n5122), .ck(clk), .q(
        \cache_data[13][45] ) );
  dp_1 \cache_data_reg[13][77]  ( .ip(n5090), .ck(clk), .q(
        \cache_data[13][77] ) );
  dp_1 \cache_data_reg[13][109]  ( .ip(n5058), .ck(clk), .q(
        \cache_data[13][109] ) );
  dp_1 \cache_data_reg[14][13]  ( .ip(n5026), .ck(clk), .q(
        \cache_data[14][13] ) );
  dp_1 \cache_data_reg[14][45]  ( .ip(n4994), .ck(clk), .q(
        \cache_data[14][45] ) );
  dp_1 \cache_data_reg[14][77]  ( .ip(n4962), .ck(clk), .q(
        \cache_data[14][77] ) );
  dp_1 \cache_data_reg[14][109]  ( .ip(n4930), .ck(clk), .q(
        \cache_data[14][109] ) );
  dp_1 \cache_data_reg[15][13]  ( .ip(n4898), .ck(clk), .q(
        \cache_data[15][13] ) );
  dp_1 \cache_data_reg[15][45]  ( .ip(n4866), .ck(clk), .q(
        \cache_data[15][45] ) );
  dp_1 \cache_data_reg[15][77]  ( .ip(n4834), .ck(clk), .q(
        \cache_data[15][77] ) );
  dp_1 \cache_data_reg[15][109]  ( .ip(n4802), .ck(clk), .q(
        \cache_data[15][109] ) );
  dp_1 \iCache_data_wr_reg[14]  ( .ip(n6849), .ck(clk), .q(iCache_data_wr[14])
         );
  dp_1 \cache_data_reg[0][14]  ( .ip(n6817), .ck(clk), .q(\cache_data[0][14] )
         );
  dp_1 \cache_data_reg[0][46]  ( .ip(n6785), .ck(clk), .q(\cache_data[0][46] )
         );
  dp_1 \cache_data_reg[0][78]  ( .ip(n6753), .ck(clk), .q(\cache_data[0][78] )
         );
  dp_1 \cache_data_reg[0][110]  ( .ip(n6721), .ck(clk), .q(
        \cache_data[0][110] ) );
  dp_1 \cache_data_reg[1][14]  ( .ip(n6689), .ck(clk), .q(\cache_data[1][14] )
         );
  dp_1 \cache_data_reg[1][46]  ( .ip(n6657), .ck(clk), .q(\cache_data[1][46] )
         );
  dp_1 \cache_data_reg[1][78]  ( .ip(n6625), .ck(clk), .q(\cache_data[1][78] )
         );
  dp_1 \cache_data_reg[1][110]  ( .ip(n6593), .ck(clk), .q(
        \cache_data[1][110] ) );
  dp_1 \cache_data_reg[2][14]  ( .ip(n6561), .ck(clk), .q(\cache_data[2][14] )
         );
  dp_1 \cache_data_reg[2][46]  ( .ip(n6529), .ck(clk), .q(\cache_data[2][46] )
         );
  dp_1 \cache_data_reg[2][78]  ( .ip(n6497), .ck(clk), .q(\cache_data[2][78] )
         );
  dp_1 \cache_data_reg[2][110]  ( .ip(n6465), .ck(clk), .q(
        \cache_data[2][110] ) );
  dp_1 \cache_data_reg[3][14]  ( .ip(n6433), .ck(clk), .q(\cache_data[3][14] )
         );
  dp_1 \cache_data_reg[3][46]  ( .ip(n6401), .ck(clk), .q(\cache_data[3][46] )
         );
  dp_1 \cache_data_reg[3][78]  ( .ip(n6369), .ck(clk), .q(\cache_data[3][78] )
         );
  dp_1 \cache_data_reg[3][110]  ( .ip(n6337), .ck(clk), .q(
        \cache_data[3][110] ) );
  dp_1 \cache_data_reg[4][14]  ( .ip(n6305), .ck(clk), .q(\cache_data[4][14] )
         );
  dp_1 \cache_data_reg[4][46]  ( .ip(n6273), .ck(clk), .q(\cache_data[4][46] )
         );
  dp_1 \cache_data_reg[4][78]  ( .ip(n6241), .ck(clk), .q(\cache_data[4][78] )
         );
  dp_1 \cache_data_reg[4][110]  ( .ip(n6209), .ck(clk), .q(
        \cache_data[4][110] ) );
  dp_1 \cache_data_reg[5][14]  ( .ip(n6177), .ck(clk), .q(\cache_data[5][14] )
         );
  dp_1 \cache_data_reg[5][46]  ( .ip(n6145), .ck(clk), .q(\cache_data[5][46] )
         );
  dp_1 \cache_data_reg[5][78]  ( .ip(n6113), .ck(clk), .q(\cache_data[5][78] )
         );
  dp_1 \cache_data_reg[5][110]  ( .ip(n6081), .ck(clk), .q(
        \cache_data[5][110] ) );
  dp_1 \cache_data_reg[6][14]  ( .ip(n6049), .ck(clk), .q(\cache_data[6][14] )
         );
  dp_1 \cache_data_reg[6][46]  ( .ip(n6017), .ck(clk), .q(\cache_data[6][46] )
         );
  dp_1 \cache_data_reg[6][78]  ( .ip(n5985), .ck(clk), .q(\cache_data[6][78] )
         );
  dp_1 \cache_data_reg[6][110]  ( .ip(n5953), .ck(clk), .q(
        \cache_data[6][110] ) );
  dp_1 \cache_data_reg[7][14]  ( .ip(n5921), .ck(clk), .q(\cache_data[7][14] )
         );
  dp_1 \cache_data_reg[7][46]  ( .ip(n5889), .ck(clk), .q(\cache_data[7][46] )
         );
  dp_1 \cache_data_reg[7][78]  ( .ip(n5857), .ck(clk), .q(\cache_data[7][78] )
         );
  dp_1 \cache_data_reg[7][110]  ( .ip(n5825), .ck(clk), .q(
        \cache_data[7][110] ) );
  dp_1 \cache_data_reg[8][14]  ( .ip(n5793), .ck(clk), .q(\cache_data[8][14] )
         );
  dp_1 \cache_data_reg[8][46]  ( .ip(n5761), .ck(clk), .q(\cache_data[8][46] )
         );
  dp_1 \cache_data_reg[8][78]  ( .ip(n5729), .ck(clk), .q(\cache_data[8][78] )
         );
  dp_1 \cache_data_reg[8][110]  ( .ip(n5697), .ck(clk), .q(
        \cache_data[8][110] ) );
  dp_1 \cache_data_reg[9][14]  ( .ip(n5665), .ck(clk), .q(\cache_data[9][14] )
         );
  dp_1 \cache_data_reg[9][46]  ( .ip(n5633), .ck(clk), .q(\cache_data[9][46] )
         );
  dp_1 \cache_data_reg[9][78]  ( .ip(n5601), .ck(clk), .q(\cache_data[9][78] )
         );
  dp_1 \cache_data_reg[9][110]  ( .ip(n5569), .ck(clk), .q(
        \cache_data[9][110] ) );
  dp_1 \cache_data_reg[10][14]  ( .ip(n5537), .ck(clk), .q(
        \cache_data[10][14] ) );
  dp_1 \cache_data_reg[10][46]  ( .ip(n5505), .ck(clk), .q(
        \cache_data[10][46] ) );
  dp_1 \cache_data_reg[10][78]  ( .ip(n5473), .ck(clk), .q(
        \cache_data[10][78] ) );
  dp_1 \cache_data_reg[10][110]  ( .ip(n5441), .ck(clk), .q(
        \cache_data[10][110] ) );
  dp_1 \cache_data_reg[11][14]  ( .ip(n5409), .ck(clk), .q(
        \cache_data[11][14] ) );
  dp_1 \cache_data_reg[11][46]  ( .ip(n5377), .ck(clk), .q(
        \cache_data[11][46] ) );
  dp_1 \cache_data_reg[11][78]  ( .ip(n5345), .ck(clk), .q(
        \cache_data[11][78] ) );
  dp_1 \cache_data_reg[11][110]  ( .ip(n5313), .ck(clk), .q(
        \cache_data[11][110] ) );
  dp_1 \cache_data_reg[12][14]  ( .ip(n5281), .ck(clk), .q(
        \cache_data[12][14] ) );
  dp_1 \cache_data_reg[12][46]  ( .ip(n5249), .ck(clk), .q(
        \cache_data[12][46] ) );
  dp_1 \cache_data_reg[12][78]  ( .ip(n5217), .ck(clk), .q(
        \cache_data[12][78] ) );
  dp_1 \cache_data_reg[12][110]  ( .ip(n5185), .ck(clk), .q(
        \cache_data[12][110] ) );
  dp_1 \cache_data_reg[13][14]  ( .ip(n5153), .ck(clk), .q(
        \cache_data[13][14] ) );
  dp_1 \cache_data_reg[13][46]  ( .ip(n5121), .ck(clk), .q(
        \cache_data[13][46] ) );
  dp_1 \cache_data_reg[13][78]  ( .ip(n5089), .ck(clk), .q(
        \cache_data[13][78] ) );
  dp_1 \cache_data_reg[13][110]  ( .ip(n5057), .ck(clk), .q(
        \cache_data[13][110] ) );
  dp_1 \cache_data_reg[14][14]  ( .ip(n5025), .ck(clk), .q(
        \cache_data[14][14] ) );
  dp_1 \cache_data_reg[14][46]  ( .ip(n4993), .ck(clk), .q(
        \cache_data[14][46] ) );
  dp_1 \cache_data_reg[14][78]  ( .ip(n4961), .ck(clk), .q(
        \cache_data[14][78] ) );
  dp_1 \cache_data_reg[14][110]  ( .ip(n4929), .ck(clk), .q(
        \cache_data[14][110] ) );
  dp_1 \cache_data_reg[15][14]  ( .ip(n4897), .ck(clk), .q(
        \cache_data[15][14] ) );
  dp_1 \cache_data_reg[15][46]  ( .ip(n4865), .ck(clk), .q(
        \cache_data[15][46] ) );
  dp_1 \cache_data_reg[15][78]  ( .ip(n4833), .ck(clk), .q(
        \cache_data[15][78] ) );
  dp_1 \cache_data_reg[15][110]  ( .ip(n4801), .ck(clk), .q(
        \cache_data[15][110] ) );
  dp_1 \iCache_data_wr_reg[15]  ( .ip(n6848), .ck(clk), .q(iCache_data_wr[15])
         );
  dp_1 \cache_data_reg[0][15]  ( .ip(n6816), .ck(clk), .q(\cache_data[0][15] )
         );
  dp_1 \cache_data_reg[0][47]  ( .ip(n6784), .ck(clk), .q(\cache_data[0][47] )
         );
  dp_1 \cache_data_reg[0][79]  ( .ip(n6752), .ck(clk), .q(\cache_data[0][79] )
         );
  dp_1 \cache_data_reg[0][111]  ( .ip(n6720), .ck(clk), .q(
        \cache_data[0][111] ) );
  dp_1 \cache_data_reg[1][15]  ( .ip(n6688), .ck(clk), .q(\cache_data[1][15] )
         );
  dp_1 \cache_data_reg[1][47]  ( .ip(n6656), .ck(clk), .q(\cache_data[1][47] )
         );
  dp_1 \cache_data_reg[1][79]  ( .ip(n6624), .ck(clk), .q(\cache_data[1][79] )
         );
  dp_1 \cache_data_reg[1][111]  ( .ip(n6592), .ck(clk), .q(
        \cache_data[1][111] ) );
  dp_1 \cache_data_reg[2][15]  ( .ip(n6560), .ck(clk), .q(\cache_data[2][15] )
         );
  dp_1 \cache_data_reg[2][47]  ( .ip(n6528), .ck(clk), .q(\cache_data[2][47] )
         );
  dp_1 \cache_data_reg[2][79]  ( .ip(n6496), .ck(clk), .q(\cache_data[2][79] )
         );
  dp_1 \cache_data_reg[2][111]  ( .ip(n6464), .ck(clk), .q(
        \cache_data[2][111] ) );
  dp_1 \cache_data_reg[3][15]  ( .ip(n6432), .ck(clk), .q(\cache_data[3][15] )
         );
  dp_1 \cache_data_reg[3][47]  ( .ip(n6400), .ck(clk), .q(\cache_data[3][47] )
         );
  dp_1 \cache_data_reg[3][79]  ( .ip(n6368), .ck(clk), .q(\cache_data[3][79] )
         );
  dp_1 \cache_data_reg[3][111]  ( .ip(n6336), .ck(clk), .q(
        \cache_data[3][111] ) );
  dp_1 \cache_data_reg[4][15]  ( .ip(n6304), .ck(clk), .q(\cache_data[4][15] )
         );
  dp_1 \cache_data_reg[4][47]  ( .ip(n6272), .ck(clk), .q(\cache_data[4][47] )
         );
  dp_1 \cache_data_reg[4][79]  ( .ip(n6240), .ck(clk), .q(\cache_data[4][79] )
         );
  dp_1 \cache_data_reg[4][111]  ( .ip(n6208), .ck(clk), .q(
        \cache_data[4][111] ) );
  dp_1 \cache_data_reg[5][15]  ( .ip(n6176), .ck(clk), .q(\cache_data[5][15] )
         );
  dp_1 \cache_data_reg[5][47]  ( .ip(n6144), .ck(clk), .q(\cache_data[5][47] )
         );
  dp_1 \cache_data_reg[5][79]  ( .ip(n6112), .ck(clk), .q(\cache_data[5][79] )
         );
  dp_1 \cache_data_reg[5][111]  ( .ip(n6080), .ck(clk), .q(
        \cache_data[5][111] ) );
  dp_1 \cache_data_reg[6][15]  ( .ip(n6048), .ck(clk), .q(\cache_data[6][15] )
         );
  dp_1 \cache_data_reg[6][47]  ( .ip(n6016), .ck(clk), .q(\cache_data[6][47] )
         );
  dp_1 \cache_data_reg[6][79]  ( .ip(n5984), .ck(clk), .q(\cache_data[6][79] )
         );
  dp_1 \cache_data_reg[6][111]  ( .ip(n5952), .ck(clk), .q(
        \cache_data[6][111] ) );
  dp_1 \cache_data_reg[7][15]  ( .ip(n5920), .ck(clk), .q(\cache_data[7][15] )
         );
  dp_1 \cache_data_reg[7][47]  ( .ip(n5888), .ck(clk), .q(\cache_data[7][47] )
         );
  dp_1 \cache_data_reg[7][79]  ( .ip(n5856), .ck(clk), .q(\cache_data[7][79] )
         );
  dp_1 \cache_data_reg[7][111]  ( .ip(n5824), .ck(clk), .q(
        \cache_data[7][111] ) );
  dp_1 \cache_data_reg[8][15]  ( .ip(n5792), .ck(clk), .q(\cache_data[8][15] )
         );
  dp_1 \cache_data_reg[8][47]  ( .ip(n5760), .ck(clk), .q(\cache_data[8][47] )
         );
  dp_1 \cache_data_reg[8][79]  ( .ip(n5728), .ck(clk), .q(\cache_data[8][79] )
         );
  dp_1 \cache_data_reg[8][111]  ( .ip(n5696), .ck(clk), .q(
        \cache_data[8][111] ) );
  dp_1 \cache_data_reg[9][15]  ( .ip(n5664), .ck(clk), .q(\cache_data[9][15] )
         );
  dp_1 \cache_data_reg[9][47]  ( .ip(n5632), .ck(clk), .q(\cache_data[9][47] )
         );
  dp_1 \cache_data_reg[9][79]  ( .ip(n5600), .ck(clk), .q(\cache_data[9][79] )
         );
  dp_1 \cache_data_reg[9][111]  ( .ip(n5568), .ck(clk), .q(
        \cache_data[9][111] ) );
  dp_1 \cache_data_reg[10][15]  ( .ip(n5536), .ck(clk), .q(
        \cache_data[10][15] ) );
  dp_1 \cache_data_reg[10][47]  ( .ip(n5504), .ck(clk), .q(
        \cache_data[10][47] ) );
  dp_1 \cache_data_reg[10][79]  ( .ip(n5472), .ck(clk), .q(
        \cache_data[10][79] ) );
  dp_1 \cache_data_reg[10][111]  ( .ip(n5440), .ck(clk), .q(
        \cache_data[10][111] ) );
  dp_1 \cache_data_reg[11][15]  ( .ip(n5408), .ck(clk), .q(
        \cache_data[11][15] ) );
  dp_1 \cache_data_reg[11][47]  ( .ip(n5376), .ck(clk), .q(
        \cache_data[11][47] ) );
  dp_1 \cache_data_reg[11][79]  ( .ip(n5344), .ck(clk), .q(
        \cache_data[11][79] ) );
  dp_1 \cache_data_reg[11][111]  ( .ip(n5312), .ck(clk), .q(
        \cache_data[11][111] ) );
  dp_1 \cache_data_reg[12][15]  ( .ip(n5280), .ck(clk), .q(
        \cache_data[12][15] ) );
  dp_1 \cache_data_reg[12][47]  ( .ip(n5248), .ck(clk), .q(
        \cache_data[12][47] ) );
  dp_1 \cache_data_reg[12][79]  ( .ip(n5216), .ck(clk), .q(
        \cache_data[12][79] ) );
  dp_1 \cache_data_reg[12][111]  ( .ip(n5184), .ck(clk), .q(
        \cache_data[12][111] ) );
  dp_1 \cache_data_reg[13][15]  ( .ip(n5152), .ck(clk), .q(
        \cache_data[13][15] ) );
  dp_1 \cache_data_reg[13][47]  ( .ip(n5120), .ck(clk), .q(
        \cache_data[13][47] ) );
  dp_1 \cache_data_reg[13][79]  ( .ip(n5088), .ck(clk), .q(
        \cache_data[13][79] ) );
  dp_1 \cache_data_reg[13][111]  ( .ip(n5056), .ck(clk), .q(
        \cache_data[13][111] ) );
  dp_1 \cache_data_reg[14][15]  ( .ip(n5024), .ck(clk), .q(
        \cache_data[14][15] ) );
  dp_1 \cache_data_reg[14][47]  ( .ip(n4992), .ck(clk), .q(
        \cache_data[14][47] ) );
  dp_1 \cache_data_reg[14][79]  ( .ip(n4960), .ck(clk), .q(
        \cache_data[14][79] ) );
  dp_1 \cache_data_reg[14][111]  ( .ip(n4928), .ck(clk), .q(
        \cache_data[14][111] ) );
  dp_1 \cache_data_reg[15][15]  ( .ip(n4896), .ck(clk), .q(
        \cache_data[15][15] ) );
  dp_1 \cache_data_reg[15][47]  ( .ip(n4864), .ck(clk), .q(
        \cache_data[15][47] ) );
  dp_1 \cache_data_reg[15][79]  ( .ip(n4832), .ck(clk), .q(
        \cache_data[15][79] ) );
  dp_1 \cache_data_reg[15][111]  ( .ip(n4800), .ck(clk), .q(
        \cache_data[15][111] ) );
  dp_1 \iCache_data_wr_reg[16]  ( .ip(n6847), .ck(clk), .q(iCache_data_wr[16])
         );
  dp_1 \cache_data_reg[0][16]  ( .ip(n6815), .ck(clk), .q(\cache_data[0][16] )
         );
  dp_1 \cache_data_reg[0][48]  ( .ip(n6783), .ck(clk), .q(\cache_data[0][48] )
         );
  dp_1 \cache_data_reg[0][80]  ( .ip(n6751), .ck(clk), .q(\cache_data[0][80] )
         );
  dp_1 \cache_data_reg[0][112]  ( .ip(n6719), .ck(clk), .q(
        \cache_data[0][112] ) );
  dp_1 \cache_data_reg[1][16]  ( .ip(n6687), .ck(clk), .q(\cache_data[1][16] )
         );
  dp_1 \cache_data_reg[1][48]  ( .ip(n6655), .ck(clk), .q(\cache_data[1][48] )
         );
  dp_1 \cache_data_reg[1][80]  ( .ip(n6623), .ck(clk), .q(\cache_data[1][80] )
         );
  dp_1 \cache_data_reg[1][112]  ( .ip(n6591), .ck(clk), .q(
        \cache_data[1][112] ) );
  dp_1 \cache_data_reg[2][16]  ( .ip(n6559), .ck(clk), .q(\cache_data[2][16] )
         );
  dp_1 \cache_data_reg[2][48]  ( .ip(n6527), .ck(clk), .q(\cache_data[2][48] )
         );
  dp_1 \cache_data_reg[2][80]  ( .ip(n6495), .ck(clk), .q(\cache_data[2][80] )
         );
  dp_1 \cache_data_reg[2][112]  ( .ip(n6463), .ck(clk), .q(
        \cache_data[2][112] ) );
  dp_1 \cache_data_reg[3][16]  ( .ip(n6431), .ck(clk), .q(\cache_data[3][16] )
         );
  dp_1 \cache_data_reg[3][48]  ( .ip(n6399), .ck(clk), .q(\cache_data[3][48] )
         );
  dp_1 \cache_data_reg[3][80]  ( .ip(n6367), .ck(clk), .q(\cache_data[3][80] )
         );
  dp_1 \cache_data_reg[3][112]  ( .ip(n6335), .ck(clk), .q(
        \cache_data[3][112] ) );
  dp_1 \cache_data_reg[4][16]  ( .ip(n6303), .ck(clk), .q(\cache_data[4][16] )
         );
  dp_1 \cache_data_reg[4][48]  ( .ip(n6271), .ck(clk), .q(\cache_data[4][48] )
         );
  dp_1 \cache_data_reg[4][80]  ( .ip(n6239), .ck(clk), .q(\cache_data[4][80] )
         );
  dp_1 \cache_data_reg[4][112]  ( .ip(n6207), .ck(clk), .q(
        \cache_data[4][112] ) );
  dp_1 \cache_data_reg[5][16]  ( .ip(n6175), .ck(clk), .q(\cache_data[5][16] )
         );
  dp_1 \cache_data_reg[5][48]  ( .ip(n6143), .ck(clk), .q(\cache_data[5][48] )
         );
  dp_1 \cache_data_reg[5][80]  ( .ip(n6111), .ck(clk), .q(\cache_data[5][80] )
         );
  dp_1 \cache_data_reg[5][112]  ( .ip(n6079), .ck(clk), .q(
        \cache_data[5][112] ) );
  dp_1 \cache_data_reg[6][16]  ( .ip(n6047), .ck(clk), .q(\cache_data[6][16] )
         );
  dp_1 \cache_data_reg[6][48]  ( .ip(n6015), .ck(clk), .q(\cache_data[6][48] )
         );
  dp_1 \cache_data_reg[6][80]  ( .ip(n5983), .ck(clk), .q(\cache_data[6][80] )
         );
  dp_1 \cache_data_reg[6][112]  ( .ip(n5951), .ck(clk), .q(
        \cache_data[6][112] ) );
  dp_1 \cache_data_reg[7][16]  ( .ip(n5919), .ck(clk), .q(\cache_data[7][16] )
         );
  dp_1 \cache_data_reg[7][48]  ( .ip(n5887), .ck(clk), .q(\cache_data[7][48] )
         );
  dp_1 \cache_data_reg[7][80]  ( .ip(n5855), .ck(clk), .q(\cache_data[7][80] )
         );
  dp_1 \cache_data_reg[7][112]  ( .ip(n5823), .ck(clk), .q(
        \cache_data[7][112] ) );
  dp_1 \cache_data_reg[8][16]  ( .ip(n5791), .ck(clk), .q(\cache_data[8][16] )
         );
  dp_1 \cache_data_reg[8][48]  ( .ip(n5759), .ck(clk), .q(\cache_data[8][48] )
         );
  dp_1 \cache_data_reg[8][80]  ( .ip(n5727), .ck(clk), .q(\cache_data[8][80] )
         );
  dp_1 \cache_data_reg[8][112]  ( .ip(n5695), .ck(clk), .q(
        \cache_data[8][112] ) );
  dp_1 \cache_data_reg[9][16]  ( .ip(n5663), .ck(clk), .q(\cache_data[9][16] )
         );
  dp_1 \cache_data_reg[9][48]  ( .ip(n5631), .ck(clk), .q(\cache_data[9][48] )
         );
  dp_1 \cache_data_reg[9][80]  ( .ip(n5599), .ck(clk), .q(\cache_data[9][80] )
         );
  dp_1 \cache_data_reg[9][112]  ( .ip(n5567), .ck(clk), .q(
        \cache_data[9][112] ) );
  dp_1 \cache_data_reg[10][16]  ( .ip(n5535), .ck(clk), .q(
        \cache_data[10][16] ) );
  dp_1 \cache_data_reg[10][48]  ( .ip(n5503), .ck(clk), .q(
        \cache_data[10][48] ) );
  dp_1 \cache_data_reg[10][80]  ( .ip(n5471), .ck(clk), .q(
        \cache_data[10][80] ) );
  dp_1 \cache_data_reg[10][112]  ( .ip(n5439), .ck(clk), .q(
        \cache_data[10][112] ) );
  dp_1 \cache_data_reg[11][16]  ( .ip(n5407), .ck(clk), .q(
        \cache_data[11][16] ) );
  dp_1 \cache_data_reg[11][48]  ( .ip(n5375), .ck(clk), .q(
        \cache_data[11][48] ) );
  dp_1 \cache_data_reg[11][80]  ( .ip(n5343), .ck(clk), .q(
        \cache_data[11][80] ) );
  dp_1 \cache_data_reg[11][112]  ( .ip(n5311), .ck(clk), .q(
        \cache_data[11][112] ) );
  dp_1 \cache_data_reg[12][16]  ( .ip(n5279), .ck(clk), .q(
        \cache_data[12][16] ) );
  dp_1 \cache_data_reg[12][48]  ( .ip(n5247), .ck(clk), .q(
        \cache_data[12][48] ) );
  dp_1 \cache_data_reg[12][80]  ( .ip(n5215), .ck(clk), .q(
        \cache_data[12][80] ) );
  dp_1 \cache_data_reg[12][112]  ( .ip(n5183), .ck(clk), .q(
        \cache_data[12][112] ) );
  dp_1 \cache_data_reg[13][16]  ( .ip(n5151), .ck(clk), .q(
        \cache_data[13][16] ) );
  dp_1 \cache_data_reg[13][48]  ( .ip(n5119), .ck(clk), .q(
        \cache_data[13][48] ) );
  dp_1 \cache_data_reg[13][80]  ( .ip(n5087), .ck(clk), .q(
        \cache_data[13][80] ) );
  dp_1 \cache_data_reg[13][112]  ( .ip(n5055), .ck(clk), .q(
        \cache_data[13][112] ) );
  dp_1 \cache_data_reg[14][16]  ( .ip(n5023), .ck(clk), .q(
        \cache_data[14][16] ) );
  dp_1 \cache_data_reg[14][48]  ( .ip(n4991), .ck(clk), .q(
        \cache_data[14][48] ) );
  dp_1 \cache_data_reg[14][80]  ( .ip(n4959), .ck(clk), .q(
        \cache_data[14][80] ) );
  dp_1 \cache_data_reg[14][112]  ( .ip(n4927), .ck(clk), .q(
        \cache_data[14][112] ) );
  dp_1 \cache_data_reg[15][16]  ( .ip(n4895), .ck(clk), .q(
        \cache_data[15][16] ) );
  dp_1 \cache_data_reg[15][48]  ( .ip(n4863), .ck(clk), .q(
        \cache_data[15][48] ) );
  dp_1 \cache_data_reg[15][80]  ( .ip(n4831), .ck(clk), .q(
        \cache_data[15][80] ) );
  dp_1 \cache_data_reg[15][112]  ( .ip(n4799), .ck(clk), .q(
        \cache_data[15][112] ) );
  dp_1 \iCache_data_wr_reg[17]  ( .ip(n6846), .ck(clk), .q(iCache_data_wr[17])
         );
  dp_1 \cache_data_reg[0][17]  ( .ip(n6814), .ck(clk), .q(\cache_data[0][17] )
         );
  dp_1 \cache_data_reg[0][49]  ( .ip(n6782), .ck(clk), .q(\cache_data[0][49] )
         );
  dp_1 \cache_data_reg[0][81]  ( .ip(n6750), .ck(clk), .q(\cache_data[0][81] )
         );
  dp_1 \cache_data_reg[0][113]  ( .ip(n6718), .ck(clk), .q(
        \cache_data[0][113] ) );
  dp_1 \cache_data_reg[1][17]  ( .ip(n6686), .ck(clk), .q(\cache_data[1][17] )
         );
  dp_1 \cache_data_reg[1][49]  ( .ip(n6654), .ck(clk), .q(\cache_data[1][49] )
         );
  dp_1 \cache_data_reg[1][81]  ( .ip(n6622), .ck(clk), .q(\cache_data[1][81] )
         );
  dp_1 \cache_data_reg[1][113]  ( .ip(n6590), .ck(clk), .q(
        \cache_data[1][113] ) );
  dp_1 \cache_data_reg[2][17]  ( .ip(n6558), .ck(clk), .q(\cache_data[2][17] )
         );
  dp_1 \cache_data_reg[2][49]  ( .ip(n6526), .ck(clk), .q(\cache_data[2][49] )
         );
  dp_1 \cache_data_reg[2][81]  ( .ip(n6494), .ck(clk), .q(\cache_data[2][81] )
         );
  dp_1 \cache_data_reg[2][113]  ( .ip(n6462), .ck(clk), .q(
        \cache_data[2][113] ) );
  dp_1 \cache_data_reg[3][17]  ( .ip(n6430), .ck(clk), .q(\cache_data[3][17] )
         );
  dp_1 \cache_data_reg[3][49]  ( .ip(n6398), .ck(clk), .q(\cache_data[3][49] )
         );
  dp_1 \cache_data_reg[3][81]  ( .ip(n6366), .ck(clk), .q(\cache_data[3][81] )
         );
  dp_1 \cache_data_reg[3][113]  ( .ip(n6334), .ck(clk), .q(
        \cache_data[3][113] ) );
  dp_1 \cache_data_reg[4][17]  ( .ip(n6302), .ck(clk), .q(\cache_data[4][17] )
         );
  dp_1 \cache_data_reg[4][49]  ( .ip(n6270), .ck(clk), .q(\cache_data[4][49] )
         );
  dp_1 \cache_data_reg[4][81]  ( .ip(n6238), .ck(clk), .q(\cache_data[4][81] )
         );
  dp_1 \cache_data_reg[4][113]  ( .ip(n6206), .ck(clk), .q(
        \cache_data[4][113] ) );
  dp_1 \cache_data_reg[5][17]  ( .ip(n6174), .ck(clk), .q(\cache_data[5][17] )
         );
  dp_1 \cache_data_reg[5][49]  ( .ip(n6142), .ck(clk), .q(\cache_data[5][49] )
         );
  dp_1 \cache_data_reg[5][81]  ( .ip(n6110), .ck(clk), .q(\cache_data[5][81] )
         );
  dp_1 \cache_data_reg[5][113]  ( .ip(n6078), .ck(clk), .q(
        \cache_data[5][113] ) );
  dp_1 \cache_data_reg[6][17]  ( .ip(n6046), .ck(clk), .q(\cache_data[6][17] )
         );
  dp_1 \cache_data_reg[6][49]  ( .ip(n6014), .ck(clk), .q(\cache_data[6][49] )
         );
  dp_1 \cache_data_reg[6][81]  ( .ip(n5982), .ck(clk), .q(\cache_data[6][81] )
         );
  dp_1 \cache_data_reg[6][113]  ( .ip(n5950), .ck(clk), .q(
        \cache_data[6][113] ) );
  dp_1 \cache_data_reg[7][17]  ( .ip(n5918), .ck(clk), .q(\cache_data[7][17] )
         );
  dp_1 \cache_data_reg[7][49]  ( .ip(n5886), .ck(clk), .q(\cache_data[7][49] )
         );
  dp_1 \cache_data_reg[7][81]  ( .ip(n5854), .ck(clk), .q(\cache_data[7][81] )
         );
  dp_1 \cache_data_reg[7][113]  ( .ip(n5822), .ck(clk), .q(
        \cache_data[7][113] ) );
  dp_1 \cache_data_reg[8][17]  ( .ip(n5790), .ck(clk), .q(\cache_data[8][17] )
         );
  dp_1 \cache_data_reg[8][49]  ( .ip(n5758), .ck(clk), .q(\cache_data[8][49] )
         );
  dp_1 \cache_data_reg[8][81]  ( .ip(n5726), .ck(clk), .q(\cache_data[8][81] )
         );
  dp_1 \cache_data_reg[8][113]  ( .ip(n5694), .ck(clk), .q(
        \cache_data[8][113] ) );
  dp_1 \cache_data_reg[9][17]  ( .ip(n5662), .ck(clk), .q(\cache_data[9][17] )
         );
  dp_1 \cache_data_reg[9][49]  ( .ip(n5630), .ck(clk), .q(\cache_data[9][49] )
         );
  dp_1 \cache_data_reg[9][81]  ( .ip(n5598), .ck(clk), .q(\cache_data[9][81] )
         );
  dp_1 \cache_data_reg[9][113]  ( .ip(n5566), .ck(clk), .q(
        \cache_data[9][113] ) );
  dp_1 \cache_data_reg[10][17]  ( .ip(n5534), .ck(clk), .q(
        \cache_data[10][17] ) );
  dp_1 \cache_data_reg[10][49]  ( .ip(n5502), .ck(clk), .q(
        \cache_data[10][49] ) );
  dp_1 \cache_data_reg[10][81]  ( .ip(n5470), .ck(clk), .q(
        \cache_data[10][81] ) );
  dp_1 \cache_data_reg[10][113]  ( .ip(n5438), .ck(clk), .q(
        \cache_data[10][113] ) );
  dp_1 \cache_data_reg[11][17]  ( .ip(n5406), .ck(clk), .q(
        \cache_data[11][17] ) );
  dp_1 \cache_data_reg[11][49]  ( .ip(n5374), .ck(clk), .q(
        \cache_data[11][49] ) );
  dp_1 \cache_data_reg[11][81]  ( .ip(n5342), .ck(clk), .q(
        \cache_data[11][81] ) );
  dp_1 \cache_data_reg[11][113]  ( .ip(n5310), .ck(clk), .q(
        \cache_data[11][113] ) );
  dp_1 \cache_data_reg[12][17]  ( .ip(n5278), .ck(clk), .q(
        \cache_data[12][17] ) );
  dp_1 \cache_data_reg[12][49]  ( .ip(n5246), .ck(clk), .q(
        \cache_data[12][49] ) );
  dp_1 \cache_data_reg[12][81]  ( .ip(n5214), .ck(clk), .q(
        \cache_data[12][81] ) );
  dp_1 \cache_data_reg[12][113]  ( .ip(n5182), .ck(clk), .q(
        \cache_data[12][113] ) );
  dp_1 \cache_data_reg[13][17]  ( .ip(n5150), .ck(clk), .q(
        \cache_data[13][17] ) );
  dp_1 \cache_data_reg[13][49]  ( .ip(n5118), .ck(clk), .q(
        \cache_data[13][49] ) );
  dp_1 \cache_data_reg[13][81]  ( .ip(n5086), .ck(clk), .q(
        \cache_data[13][81] ) );
  dp_1 \cache_data_reg[13][113]  ( .ip(n5054), .ck(clk), .q(
        \cache_data[13][113] ) );
  dp_1 \cache_data_reg[14][17]  ( .ip(n5022), .ck(clk), .q(
        \cache_data[14][17] ) );
  dp_1 \cache_data_reg[14][49]  ( .ip(n4990), .ck(clk), .q(
        \cache_data[14][49] ) );
  dp_1 \cache_data_reg[14][81]  ( .ip(n4958), .ck(clk), .q(
        \cache_data[14][81] ) );
  dp_1 \cache_data_reg[14][113]  ( .ip(n4926), .ck(clk), .q(
        \cache_data[14][113] ) );
  dp_1 \cache_data_reg[15][17]  ( .ip(n4894), .ck(clk), .q(
        \cache_data[15][17] ) );
  dp_1 \cache_data_reg[15][49]  ( .ip(n4862), .ck(clk), .q(
        \cache_data[15][49] ) );
  dp_1 \cache_data_reg[15][81]  ( .ip(n4830), .ck(clk), .q(
        \cache_data[15][81] ) );
  dp_1 \cache_data_reg[15][113]  ( .ip(n4798), .ck(clk), .q(
        \cache_data[15][113] ) );
  dp_1 \iCache_data_wr_reg[18]  ( .ip(n6845), .ck(clk), .q(iCache_data_wr[18])
         );
  dp_1 \cache_data_reg[0][18]  ( .ip(n6813), .ck(clk), .q(\cache_data[0][18] )
         );
  dp_1 \cache_data_reg[0][50]  ( .ip(n6781), .ck(clk), .q(\cache_data[0][50] )
         );
  dp_1 \cache_data_reg[0][82]  ( .ip(n6749), .ck(clk), .q(\cache_data[0][82] )
         );
  dp_1 \cache_data_reg[0][114]  ( .ip(n6717), .ck(clk), .q(
        \cache_data[0][114] ) );
  dp_1 \cache_data_reg[1][18]  ( .ip(n6685), .ck(clk), .q(\cache_data[1][18] )
         );
  dp_1 \cache_data_reg[1][50]  ( .ip(n6653), .ck(clk), .q(\cache_data[1][50] )
         );
  dp_1 \cache_data_reg[1][82]  ( .ip(n6621), .ck(clk), .q(\cache_data[1][82] )
         );
  dp_1 \cache_data_reg[1][114]  ( .ip(n6589), .ck(clk), .q(
        \cache_data[1][114] ) );
  dp_1 \cache_data_reg[2][18]  ( .ip(n6557), .ck(clk), .q(\cache_data[2][18] )
         );
  dp_1 \cache_data_reg[2][50]  ( .ip(n6525), .ck(clk), .q(\cache_data[2][50] )
         );
  dp_1 \cache_data_reg[2][82]  ( .ip(n6493), .ck(clk), .q(\cache_data[2][82] )
         );
  dp_1 \cache_data_reg[2][114]  ( .ip(n6461), .ck(clk), .q(
        \cache_data[2][114] ) );
  dp_1 \cache_data_reg[3][18]  ( .ip(n6429), .ck(clk), .q(\cache_data[3][18] )
         );
  dp_1 \cache_data_reg[3][50]  ( .ip(n6397), .ck(clk), .q(\cache_data[3][50] )
         );
  dp_1 \cache_data_reg[3][82]  ( .ip(n6365), .ck(clk), .q(\cache_data[3][82] )
         );
  dp_1 \cache_data_reg[3][114]  ( .ip(n6333), .ck(clk), .q(
        \cache_data[3][114] ) );
  dp_1 \cache_data_reg[4][18]  ( .ip(n6301), .ck(clk), .q(\cache_data[4][18] )
         );
  dp_1 \cache_data_reg[4][50]  ( .ip(n6269), .ck(clk), .q(\cache_data[4][50] )
         );
  dp_1 \cache_data_reg[4][82]  ( .ip(n6237), .ck(clk), .q(\cache_data[4][82] )
         );
  dp_1 \cache_data_reg[4][114]  ( .ip(n6205), .ck(clk), .q(
        \cache_data[4][114] ) );
  dp_1 \cache_data_reg[5][18]  ( .ip(n6173), .ck(clk), .q(\cache_data[5][18] )
         );
  dp_1 \cache_data_reg[5][50]  ( .ip(n6141), .ck(clk), .q(\cache_data[5][50] )
         );
  dp_1 \cache_data_reg[5][82]  ( .ip(n6109), .ck(clk), .q(\cache_data[5][82] )
         );
  dp_1 \cache_data_reg[5][114]  ( .ip(n6077), .ck(clk), .q(
        \cache_data[5][114] ) );
  dp_1 \cache_data_reg[6][18]  ( .ip(n6045), .ck(clk), .q(\cache_data[6][18] )
         );
  dp_1 \cache_data_reg[6][50]  ( .ip(n6013), .ck(clk), .q(\cache_data[6][50] )
         );
  dp_1 \cache_data_reg[6][82]  ( .ip(n5981), .ck(clk), .q(\cache_data[6][82] )
         );
  dp_1 \cache_data_reg[6][114]  ( .ip(n5949), .ck(clk), .q(
        \cache_data[6][114] ) );
  dp_1 \cache_data_reg[7][18]  ( .ip(n5917), .ck(clk), .q(\cache_data[7][18] )
         );
  dp_1 \cache_data_reg[7][50]  ( .ip(n5885), .ck(clk), .q(\cache_data[7][50] )
         );
  dp_1 \cache_data_reg[7][82]  ( .ip(n5853), .ck(clk), .q(\cache_data[7][82] )
         );
  dp_1 \cache_data_reg[7][114]  ( .ip(n5821), .ck(clk), .q(
        \cache_data[7][114] ) );
  dp_1 \cache_data_reg[8][18]  ( .ip(n5789), .ck(clk), .q(\cache_data[8][18] )
         );
  dp_1 \cache_data_reg[8][50]  ( .ip(n5757), .ck(clk), .q(\cache_data[8][50] )
         );
  dp_1 \cache_data_reg[8][82]  ( .ip(n5725), .ck(clk), .q(\cache_data[8][82] )
         );
  dp_1 \cache_data_reg[8][114]  ( .ip(n5693), .ck(clk), .q(
        \cache_data[8][114] ) );
  dp_1 \cache_data_reg[9][18]  ( .ip(n5661), .ck(clk), .q(\cache_data[9][18] )
         );
  dp_1 \cache_data_reg[9][50]  ( .ip(n5629), .ck(clk), .q(\cache_data[9][50] )
         );
  dp_1 \cache_data_reg[9][82]  ( .ip(n5597), .ck(clk), .q(\cache_data[9][82] )
         );
  dp_1 \cache_data_reg[9][114]  ( .ip(n5565), .ck(clk), .q(
        \cache_data[9][114] ) );
  dp_1 \cache_data_reg[10][18]  ( .ip(n5533), .ck(clk), .q(
        \cache_data[10][18] ) );
  dp_1 \cache_data_reg[10][50]  ( .ip(n5501), .ck(clk), .q(
        \cache_data[10][50] ) );
  dp_1 \cache_data_reg[10][82]  ( .ip(n5469), .ck(clk), .q(
        \cache_data[10][82] ) );
  dp_1 \cache_data_reg[10][114]  ( .ip(n5437), .ck(clk), .q(
        \cache_data[10][114] ) );
  dp_1 \cache_data_reg[11][18]  ( .ip(n5405), .ck(clk), .q(
        \cache_data[11][18] ) );
  dp_1 \cache_data_reg[11][50]  ( .ip(n5373), .ck(clk), .q(
        \cache_data[11][50] ) );
  dp_1 \cache_data_reg[11][82]  ( .ip(n5341), .ck(clk), .q(
        \cache_data[11][82] ) );
  dp_1 \cache_data_reg[11][114]  ( .ip(n5309), .ck(clk), .q(
        \cache_data[11][114] ) );
  dp_1 \cache_data_reg[12][18]  ( .ip(n5277), .ck(clk), .q(
        \cache_data[12][18] ) );
  dp_1 \cache_data_reg[12][50]  ( .ip(n5245), .ck(clk), .q(
        \cache_data[12][50] ) );
  dp_1 \cache_data_reg[12][82]  ( .ip(n5213), .ck(clk), .q(
        \cache_data[12][82] ) );
  dp_1 \cache_data_reg[12][114]  ( .ip(n5181), .ck(clk), .q(
        \cache_data[12][114] ) );
  dp_1 \cache_data_reg[13][18]  ( .ip(n5149), .ck(clk), .q(
        \cache_data[13][18] ) );
  dp_1 \cache_data_reg[13][50]  ( .ip(n5117), .ck(clk), .q(
        \cache_data[13][50] ) );
  dp_1 \cache_data_reg[13][82]  ( .ip(n5085), .ck(clk), .q(
        \cache_data[13][82] ) );
  dp_1 \cache_data_reg[13][114]  ( .ip(n5053), .ck(clk), .q(
        \cache_data[13][114] ) );
  dp_1 \cache_data_reg[14][18]  ( .ip(n5021), .ck(clk), .q(
        \cache_data[14][18] ) );
  dp_1 \cache_data_reg[14][50]  ( .ip(n4989), .ck(clk), .q(
        \cache_data[14][50] ) );
  dp_1 \cache_data_reg[14][82]  ( .ip(n4957), .ck(clk), .q(
        \cache_data[14][82] ) );
  dp_1 \cache_data_reg[14][114]  ( .ip(n4925), .ck(clk), .q(
        \cache_data[14][114] ) );
  dp_1 \cache_data_reg[15][18]  ( .ip(n4893), .ck(clk), .q(
        \cache_data[15][18] ) );
  dp_1 \cache_data_reg[15][50]  ( .ip(n4861), .ck(clk), .q(
        \cache_data[15][50] ) );
  dp_1 \cache_data_reg[15][82]  ( .ip(n4829), .ck(clk), .q(
        \cache_data[15][82] ) );
  dp_1 \cache_data_reg[15][114]  ( .ip(n4797), .ck(clk), .q(
        \cache_data[15][114] ) );
  dp_1 \iCache_data_wr_reg[19]  ( .ip(n6844), .ck(clk), .q(iCache_data_wr[19])
         );
  dp_1 \cache_data_reg[0][19]  ( .ip(n6812), .ck(clk), .q(\cache_data[0][19] )
         );
  dp_1 \cache_data_reg[0][51]  ( .ip(n6780), .ck(clk), .q(\cache_data[0][51] )
         );
  dp_1 \cache_data_reg[0][83]  ( .ip(n6748), .ck(clk), .q(\cache_data[0][83] )
         );
  dp_1 \cache_data_reg[0][115]  ( .ip(n6716), .ck(clk), .q(
        \cache_data[0][115] ) );
  dp_1 \cache_data_reg[1][19]  ( .ip(n6684), .ck(clk), .q(\cache_data[1][19] )
         );
  dp_1 \cache_data_reg[1][51]  ( .ip(n6652), .ck(clk), .q(\cache_data[1][51] )
         );
  dp_1 \cache_data_reg[1][83]  ( .ip(n6620), .ck(clk), .q(\cache_data[1][83] )
         );
  dp_1 \cache_data_reg[1][115]  ( .ip(n6588), .ck(clk), .q(
        \cache_data[1][115] ) );
  dp_1 \cache_data_reg[2][19]  ( .ip(n6556), .ck(clk), .q(\cache_data[2][19] )
         );
  dp_1 \cache_data_reg[2][51]  ( .ip(n6524), .ck(clk), .q(\cache_data[2][51] )
         );
  dp_1 \cache_data_reg[2][83]  ( .ip(n6492), .ck(clk), .q(\cache_data[2][83] )
         );
  dp_1 \cache_data_reg[2][115]  ( .ip(n6460), .ck(clk), .q(
        \cache_data[2][115] ) );
  dp_1 \cache_data_reg[3][19]  ( .ip(n6428), .ck(clk), .q(\cache_data[3][19] )
         );
  dp_1 \cache_data_reg[3][51]  ( .ip(n6396), .ck(clk), .q(\cache_data[3][51] )
         );
  dp_1 \cache_data_reg[3][83]  ( .ip(n6364), .ck(clk), .q(\cache_data[3][83] )
         );
  dp_1 \cache_data_reg[3][115]  ( .ip(n6332), .ck(clk), .q(
        \cache_data[3][115] ) );
  dp_1 \cache_data_reg[4][19]  ( .ip(n6300), .ck(clk), .q(\cache_data[4][19] )
         );
  dp_1 \cache_data_reg[4][51]  ( .ip(n6268), .ck(clk), .q(\cache_data[4][51] )
         );
  dp_1 \cache_data_reg[4][83]  ( .ip(n6236), .ck(clk), .q(\cache_data[4][83] )
         );
  dp_1 \cache_data_reg[4][115]  ( .ip(n6204), .ck(clk), .q(
        \cache_data[4][115] ) );
  dp_1 \cache_data_reg[5][19]  ( .ip(n6172), .ck(clk), .q(\cache_data[5][19] )
         );
  dp_1 \cache_data_reg[5][51]  ( .ip(n6140), .ck(clk), .q(\cache_data[5][51] )
         );
  dp_1 \cache_data_reg[5][83]  ( .ip(n6108), .ck(clk), .q(\cache_data[5][83] )
         );
  dp_1 \cache_data_reg[5][115]  ( .ip(n6076), .ck(clk), .q(
        \cache_data[5][115] ) );
  dp_1 \cache_data_reg[6][19]  ( .ip(n6044), .ck(clk), .q(\cache_data[6][19] )
         );
  dp_1 \cache_data_reg[6][51]  ( .ip(n6012), .ck(clk), .q(\cache_data[6][51] )
         );
  dp_1 \cache_data_reg[6][83]  ( .ip(n5980), .ck(clk), .q(\cache_data[6][83] )
         );
  dp_1 \cache_data_reg[6][115]  ( .ip(n5948), .ck(clk), .q(
        \cache_data[6][115] ) );
  dp_1 \cache_data_reg[7][19]  ( .ip(n5916), .ck(clk), .q(\cache_data[7][19] )
         );
  dp_1 \cache_data_reg[7][51]  ( .ip(n5884), .ck(clk), .q(\cache_data[7][51] )
         );
  dp_1 \cache_data_reg[7][83]  ( .ip(n5852), .ck(clk), .q(\cache_data[7][83] )
         );
  dp_1 \cache_data_reg[7][115]  ( .ip(n5820), .ck(clk), .q(
        \cache_data[7][115] ) );
  dp_1 \cache_data_reg[8][19]  ( .ip(n5788), .ck(clk), .q(\cache_data[8][19] )
         );
  dp_1 \cache_data_reg[8][51]  ( .ip(n5756), .ck(clk), .q(\cache_data[8][51] )
         );
  dp_1 \cache_data_reg[8][83]  ( .ip(n5724), .ck(clk), .q(\cache_data[8][83] )
         );
  dp_1 \cache_data_reg[8][115]  ( .ip(n5692), .ck(clk), .q(
        \cache_data[8][115] ) );
  dp_1 \cache_data_reg[9][19]  ( .ip(n5660), .ck(clk), .q(\cache_data[9][19] )
         );
  dp_1 \cache_data_reg[9][51]  ( .ip(n5628), .ck(clk), .q(\cache_data[9][51] )
         );
  dp_1 \cache_data_reg[9][83]  ( .ip(n5596), .ck(clk), .q(\cache_data[9][83] )
         );
  dp_1 \cache_data_reg[9][115]  ( .ip(n5564), .ck(clk), .q(
        \cache_data[9][115] ) );
  dp_1 \cache_data_reg[10][19]  ( .ip(n5532), .ck(clk), .q(
        \cache_data[10][19] ) );
  dp_1 \cache_data_reg[10][51]  ( .ip(n5500), .ck(clk), .q(
        \cache_data[10][51] ) );
  dp_1 \cache_data_reg[10][83]  ( .ip(n5468), .ck(clk), .q(
        \cache_data[10][83] ) );
  dp_1 \cache_data_reg[10][115]  ( .ip(n5436), .ck(clk), .q(
        \cache_data[10][115] ) );
  dp_1 \cache_data_reg[11][19]  ( .ip(n5404), .ck(clk), .q(
        \cache_data[11][19] ) );
  dp_1 \cache_data_reg[11][51]  ( .ip(n5372), .ck(clk), .q(
        \cache_data[11][51] ) );
  dp_1 \cache_data_reg[11][83]  ( .ip(n5340), .ck(clk), .q(
        \cache_data[11][83] ) );
  dp_1 \cache_data_reg[11][115]  ( .ip(n5308), .ck(clk), .q(
        \cache_data[11][115] ) );
  dp_1 \cache_data_reg[12][19]  ( .ip(n5276), .ck(clk), .q(
        \cache_data[12][19] ) );
  dp_1 \cache_data_reg[12][51]  ( .ip(n5244), .ck(clk), .q(
        \cache_data[12][51] ) );
  dp_1 \cache_data_reg[12][83]  ( .ip(n5212), .ck(clk), .q(
        \cache_data[12][83] ) );
  dp_1 \cache_data_reg[12][115]  ( .ip(n5180), .ck(clk), .q(
        \cache_data[12][115] ) );
  dp_1 \cache_data_reg[13][19]  ( .ip(n5148), .ck(clk), .q(
        \cache_data[13][19] ) );
  dp_1 \cache_data_reg[13][51]  ( .ip(n5116), .ck(clk), .q(
        \cache_data[13][51] ) );
  dp_1 \cache_data_reg[13][83]  ( .ip(n5084), .ck(clk), .q(
        \cache_data[13][83] ) );
  dp_1 \cache_data_reg[13][115]  ( .ip(n5052), .ck(clk), .q(
        \cache_data[13][115] ) );
  dp_1 \cache_data_reg[14][19]  ( .ip(n5020), .ck(clk), .q(
        \cache_data[14][19] ) );
  dp_1 \cache_data_reg[14][51]  ( .ip(n4988), .ck(clk), .q(
        \cache_data[14][51] ) );
  dp_1 \cache_data_reg[14][83]  ( .ip(n4956), .ck(clk), .q(
        \cache_data[14][83] ) );
  dp_1 \cache_data_reg[14][115]  ( .ip(n4924), .ck(clk), .q(
        \cache_data[14][115] ) );
  dp_1 \cache_data_reg[15][19]  ( .ip(n4892), .ck(clk), .q(
        \cache_data[15][19] ) );
  dp_1 \cache_data_reg[15][51]  ( .ip(n4860), .ck(clk), .q(
        \cache_data[15][51] ) );
  dp_1 \cache_data_reg[15][83]  ( .ip(n4828), .ck(clk), .q(
        \cache_data[15][83] ) );
  dp_1 \cache_data_reg[15][115]  ( .ip(n4796), .ck(clk), .q(
        \cache_data[15][115] ) );
  dp_1 \iCache_data_wr_reg[20]  ( .ip(n6843), .ck(clk), .q(iCache_data_wr[20])
         );
  dp_1 \cache_data_reg[0][20]  ( .ip(n6811), .ck(clk), .q(\cache_data[0][20] )
         );
  dp_1 \cache_data_reg[0][52]  ( .ip(n6779), .ck(clk), .q(\cache_data[0][52] )
         );
  dp_1 \cache_data_reg[0][84]  ( .ip(n6747), .ck(clk), .q(\cache_data[0][84] )
         );
  dp_1 \cache_data_reg[0][116]  ( .ip(n6715), .ck(clk), .q(
        \cache_data[0][116] ) );
  dp_1 \cache_data_reg[1][20]  ( .ip(n6683), .ck(clk), .q(\cache_data[1][20] )
         );
  dp_1 \cache_data_reg[1][52]  ( .ip(n6651), .ck(clk), .q(\cache_data[1][52] )
         );
  dp_1 \cache_data_reg[1][84]  ( .ip(n6619), .ck(clk), .q(\cache_data[1][84] )
         );
  dp_1 \cache_data_reg[1][116]  ( .ip(n6587), .ck(clk), .q(
        \cache_data[1][116] ) );
  dp_1 \cache_data_reg[2][20]  ( .ip(n6555), .ck(clk), .q(\cache_data[2][20] )
         );
  dp_1 \cache_data_reg[2][52]  ( .ip(n6523), .ck(clk), .q(\cache_data[2][52] )
         );
  dp_1 \cache_data_reg[2][84]  ( .ip(n6491), .ck(clk), .q(\cache_data[2][84] )
         );
  dp_1 \cache_data_reg[2][116]  ( .ip(n6459), .ck(clk), .q(
        \cache_data[2][116] ) );
  dp_1 \cache_data_reg[3][20]  ( .ip(n6427), .ck(clk), .q(\cache_data[3][20] )
         );
  dp_1 \cache_data_reg[3][52]  ( .ip(n6395), .ck(clk), .q(\cache_data[3][52] )
         );
  dp_1 \cache_data_reg[3][84]  ( .ip(n6363), .ck(clk), .q(\cache_data[3][84] )
         );
  dp_1 \cache_data_reg[3][116]  ( .ip(n6331), .ck(clk), .q(
        \cache_data[3][116] ) );
  dp_1 \cache_data_reg[4][20]  ( .ip(n6299), .ck(clk), .q(\cache_data[4][20] )
         );
  dp_1 \cache_data_reg[4][52]  ( .ip(n6267), .ck(clk), .q(\cache_data[4][52] )
         );
  dp_1 \cache_data_reg[4][84]  ( .ip(n6235), .ck(clk), .q(\cache_data[4][84] )
         );
  dp_1 \cache_data_reg[4][116]  ( .ip(n6203), .ck(clk), .q(
        \cache_data[4][116] ) );
  dp_1 \cache_data_reg[5][20]  ( .ip(n6171), .ck(clk), .q(\cache_data[5][20] )
         );
  dp_1 \cache_data_reg[5][52]  ( .ip(n6139), .ck(clk), .q(\cache_data[5][52] )
         );
  dp_1 \cache_data_reg[5][84]  ( .ip(n6107), .ck(clk), .q(\cache_data[5][84] )
         );
  dp_1 \cache_data_reg[5][116]  ( .ip(n6075), .ck(clk), .q(
        \cache_data[5][116] ) );
  dp_1 \cache_data_reg[6][20]  ( .ip(n6043), .ck(clk), .q(\cache_data[6][20] )
         );
  dp_1 \cache_data_reg[6][52]  ( .ip(n6011), .ck(clk), .q(\cache_data[6][52] )
         );
  dp_1 \cache_data_reg[6][84]  ( .ip(n5979), .ck(clk), .q(\cache_data[6][84] )
         );
  dp_1 \cache_data_reg[6][116]  ( .ip(n5947), .ck(clk), .q(
        \cache_data[6][116] ) );
  dp_1 \cache_data_reg[7][20]  ( .ip(n5915), .ck(clk), .q(\cache_data[7][20] )
         );
  dp_1 \cache_data_reg[7][52]  ( .ip(n5883), .ck(clk), .q(\cache_data[7][52] )
         );
  dp_1 \cache_data_reg[7][84]  ( .ip(n5851), .ck(clk), .q(\cache_data[7][84] )
         );
  dp_1 \cache_data_reg[7][116]  ( .ip(n5819), .ck(clk), .q(
        \cache_data[7][116] ) );
  dp_1 \cache_data_reg[8][20]  ( .ip(n5787), .ck(clk), .q(\cache_data[8][20] )
         );
  dp_1 \cache_data_reg[8][52]  ( .ip(n5755), .ck(clk), .q(\cache_data[8][52] )
         );
  dp_1 \cache_data_reg[8][84]  ( .ip(n5723), .ck(clk), .q(\cache_data[8][84] )
         );
  dp_1 \cache_data_reg[8][116]  ( .ip(n5691), .ck(clk), .q(
        \cache_data[8][116] ) );
  dp_1 \cache_data_reg[9][20]  ( .ip(n5659), .ck(clk), .q(\cache_data[9][20] )
         );
  dp_1 \cache_data_reg[9][52]  ( .ip(n5627), .ck(clk), .q(\cache_data[9][52] )
         );
  dp_1 \cache_data_reg[9][84]  ( .ip(n5595), .ck(clk), .q(\cache_data[9][84] )
         );
  dp_1 \cache_data_reg[9][116]  ( .ip(n5563), .ck(clk), .q(
        \cache_data[9][116] ) );
  dp_1 \cache_data_reg[10][20]  ( .ip(n5531), .ck(clk), .q(
        \cache_data[10][20] ) );
  dp_1 \cache_data_reg[10][52]  ( .ip(n5499), .ck(clk), .q(
        \cache_data[10][52] ) );
  dp_1 \cache_data_reg[10][84]  ( .ip(n5467), .ck(clk), .q(
        \cache_data[10][84] ) );
  dp_1 \cache_data_reg[10][116]  ( .ip(n5435), .ck(clk), .q(
        \cache_data[10][116] ) );
  dp_1 \cache_data_reg[11][20]  ( .ip(n5403), .ck(clk), .q(
        \cache_data[11][20] ) );
  dp_1 \cache_data_reg[11][52]  ( .ip(n5371), .ck(clk), .q(
        \cache_data[11][52] ) );
  dp_1 \cache_data_reg[11][84]  ( .ip(n5339), .ck(clk), .q(
        \cache_data[11][84] ) );
  dp_1 \cache_data_reg[11][116]  ( .ip(n5307), .ck(clk), .q(
        \cache_data[11][116] ) );
  dp_1 \cache_data_reg[12][20]  ( .ip(n5275), .ck(clk), .q(
        \cache_data[12][20] ) );
  dp_1 \cache_data_reg[12][52]  ( .ip(n5243), .ck(clk), .q(
        \cache_data[12][52] ) );
  dp_1 \cache_data_reg[12][84]  ( .ip(n5211), .ck(clk), .q(
        \cache_data[12][84] ) );
  dp_1 \cache_data_reg[12][116]  ( .ip(n5179), .ck(clk), .q(
        \cache_data[12][116] ) );
  dp_1 \cache_data_reg[13][20]  ( .ip(n5147), .ck(clk), .q(
        \cache_data[13][20] ) );
  dp_1 \cache_data_reg[13][52]  ( .ip(n5115), .ck(clk), .q(
        \cache_data[13][52] ) );
  dp_1 \cache_data_reg[13][84]  ( .ip(n5083), .ck(clk), .q(
        \cache_data[13][84] ) );
  dp_1 \cache_data_reg[13][116]  ( .ip(n5051), .ck(clk), .q(
        \cache_data[13][116] ) );
  dp_1 \cache_data_reg[14][20]  ( .ip(n5019), .ck(clk), .q(
        \cache_data[14][20] ) );
  dp_1 \cache_data_reg[14][52]  ( .ip(n4987), .ck(clk), .q(
        \cache_data[14][52] ) );
  dp_1 \cache_data_reg[14][84]  ( .ip(n4955), .ck(clk), .q(
        \cache_data[14][84] ) );
  dp_1 \cache_data_reg[14][116]  ( .ip(n4923), .ck(clk), .q(
        \cache_data[14][116] ) );
  dp_1 \cache_data_reg[15][20]  ( .ip(n4891), .ck(clk), .q(
        \cache_data[15][20] ) );
  dp_1 \cache_data_reg[15][52]  ( .ip(n4859), .ck(clk), .q(
        \cache_data[15][52] ) );
  dp_1 \cache_data_reg[15][84]  ( .ip(n4827), .ck(clk), .q(
        \cache_data[15][84] ) );
  dp_1 \cache_data_reg[15][116]  ( .ip(n4795), .ck(clk), .q(
        \cache_data[15][116] ) );
  dp_1 \iCache_data_wr_reg[21]  ( .ip(n6842), .ck(clk), .q(iCache_data_wr[21])
         );
  dp_1 \cache_data_reg[0][21]  ( .ip(n6810), .ck(clk), .q(\cache_data[0][21] )
         );
  dp_1 \cache_data_reg[0][53]  ( .ip(n6778), .ck(clk), .q(\cache_data[0][53] )
         );
  dp_1 \cache_data_reg[0][85]  ( .ip(n6746), .ck(clk), .q(\cache_data[0][85] )
         );
  dp_1 \cache_data_reg[0][117]  ( .ip(n6714), .ck(clk), .q(
        \cache_data[0][117] ) );
  dp_1 \cache_data_reg[1][21]  ( .ip(n6682), .ck(clk), .q(\cache_data[1][21] )
         );
  dp_1 \cache_data_reg[1][53]  ( .ip(n6650), .ck(clk), .q(\cache_data[1][53] )
         );
  dp_1 \cache_data_reg[1][85]  ( .ip(n6618), .ck(clk), .q(\cache_data[1][85] )
         );
  dp_1 \cache_data_reg[1][117]  ( .ip(n6586), .ck(clk), .q(
        \cache_data[1][117] ) );
  dp_1 \cache_data_reg[2][21]  ( .ip(n6554), .ck(clk), .q(\cache_data[2][21] )
         );
  dp_1 \cache_data_reg[2][53]  ( .ip(n6522), .ck(clk), .q(\cache_data[2][53] )
         );
  dp_1 \cache_data_reg[2][85]  ( .ip(n6490), .ck(clk), .q(\cache_data[2][85] )
         );
  dp_1 \cache_data_reg[2][117]  ( .ip(n6458), .ck(clk), .q(
        \cache_data[2][117] ) );
  dp_1 \cache_data_reg[3][21]  ( .ip(n6426), .ck(clk), .q(\cache_data[3][21] )
         );
  dp_1 \cache_data_reg[3][53]  ( .ip(n6394), .ck(clk), .q(\cache_data[3][53] )
         );
  dp_1 \cache_data_reg[3][85]  ( .ip(n6362), .ck(clk), .q(\cache_data[3][85] )
         );
  dp_1 \cache_data_reg[3][117]  ( .ip(n6330), .ck(clk), .q(
        \cache_data[3][117] ) );
  dp_1 \cache_data_reg[4][21]  ( .ip(n6298), .ck(clk), .q(\cache_data[4][21] )
         );
  dp_1 \cache_data_reg[4][53]  ( .ip(n6266), .ck(clk), .q(\cache_data[4][53] )
         );
  dp_1 \cache_data_reg[4][85]  ( .ip(n6234), .ck(clk), .q(\cache_data[4][85] )
         );
  dp_1 \cache_data_reg[4][117]  ( .ip(n6202), .ck(clk), .q(
        \cache_data[4][117] ) );
  dp_1 \cache_data_reg[5][21]  ( .ip(n6170), .ck(clk), .q(\cache_data[5][21] )
         );
  dp_1 \cache_data_reg[5][53]  ( .ip(n6138), .ck(clk), .q(\cache_data[5][53] )
         );
  dp_1 \cache_data_reg[5][85]  ( .ip(n6106), .ck(clk), .q(\cache_data[5][85] )
         );
  dp_1 \cache_data_reg[5][117]  ( .ip(n6074), .ck(clk), .q(
        \cache_data[5][117] ) );
  dp_1 \cache_data_reg[6][21]  ( .ip(n6042), .ck(clk), .q(\cache_data[6][21] )
         );
  dp_1 \cache_data_reg[6][53]  ( .ip(n6010), .ck(clk), .q(\cache_data[6][53] )
         );
  dp_1 \cache_data_reg[6][85]  ( .ip(n5978), .ck(clk), .q(\cache_data[6][85] )
         );
  dp_1 \cache_data_reg[6][117]  ( .ip(n5946), .ck(clk), .q(
        \cache_data[6][117] ) );
  dp_1 \cache_data_reg[7][21]  ( .ip(n5914), .ck(clk), .q(\cache_data[7][21] )
         );
  dp_1 \cache_data_reg[7][53]  ( .ip(n5882), .ck(clk), .q(\cache_data[7][53] )
         );
  dp_1 \cache_data_reg[7][85]  ( .ip(n5850), .ck(clk), .q(\cache_data[7][85] )
         );
  dp_1 \cache_data_reg[7][117]  ( .ip(n5818), .ck(clk), .q(
        \cache_data[7][117] ) );
  dp_1 \cache_data_reg[8][21]  ( .ip(n5786), .ck(clk), .q(\cache_data[8][21] )
         );
  dp_1 \cache_data_reg[8][53]  ( .ip(n5754), .ck(clk), .q(\cache_data[8][53] )
         );
  dp_1 \cache_data_reg[8][85]  ( .ip(n5722), .ck(clk), .q(\cache_data[8][85] )
         );
  dp_1 \cache_data_reg[8][117]  ( .ip(n5690), .ck(clk), .q(
        \cache_data[8][117] ) );
  dp_1 \cache_data_reg[9][21]  ( .ip(n5658), .ck(clk), .q(\cache_data[9][21] )
         );
  dp_1 \cache_data_reg[9][53]  ( .ip(n5626), .ck(clk), .q(\cache_data[9][53] )
         );
  dp_1 \cache_data_reg[9][85]  ( .ip(n5594), .ck(clk), .q(\cache_data[9][85] )
         );
  dp_1 \cache_data_reg[9][117]  ( .ip(n5562), .ck(clk), .q(
        \cache_data[9][117] ) );
  dp_1 \cache_data_reg[10][21]  ( .ip(n5530), .ck(clk), .q(
        \cache_data[10][21] ) );
  dp_1 \cache_data_reg[10][53]  ( .ip(n5498), .ck(clk), .q(
        \cache_data[10][53] ) );
  dp_1 \cache_data_reg[10][85]  ( .ip(n5466), .ck(clk), .q(
        \cache_data[10][85] ) );
  dp_1 \cache_data_reg[10][117]  ( .ip(n5434), .ck(clk), .q(
        \cache_data[10][117] ) );
  dp_1 \cache_data_reg[11][21]  ( .ip(n5402), .ck(clk), .q(
        \cache_data[11][21] ) );
  dp_1 \cache_data_reg[11][53]  ( .ip(n5370), .ck(clk), .q(
        \cache_data[11][53] ) );
  dp_1 \cache_data_reg[11][85]  ( .ip(n5338), .ck(clk), .q(
        \cache_data[11][85] ) );
  dp_1 \cache_data_reg[11][117]  ( .ip(n5306), .ck(clk), .q(
        \cache_data[11][117] ) );
  dp_1 \cache_data_reg[12][21]  ( .ip(n5274), .ck(clk), .q(
        \cache_data[12][21] ) );
  dp_1 \cache_data_reg[12][53]  ( .ip(n5242), .ck(clk), .q(
        \cache_data[12][53] ) );
  dp_1 \cache_data_reg[12][85]  ( .ip(n5210), .ck(clk), .q(
        \cache_data[12][85] ) );
  dp_1 \cache_data_reg[12][117]  ( .ip(n5178), .ck(clk), .q(
        \cache_data[12][117] ) );
  dp_1 \cache_data_reg[13][21]  ( .ip(n5146), .ck(clk), .q(
        \cache_data[13][21] ) );
  dp_1 \cache_data_reg[13][53]  ( .ip(n5114), .ck(clk), .q(
        \cache_data[13][53] ) );
  dp_1 \cache_data_reg[13][85]  ( .ip(n5082), .ck(clk), .q(
        \cache_data[13][85] ) );
  dp_1 \cache_data_reg[13][117]  ( .ip(n5050), .ck(clk), .q(
        \cache_data[13][117] ) );
  dp_1 \cache_data_reg[14][21]  ( .ip(n5018), .ck(clk), .q(
        \cache_data[14][21] ) );
  dp_1 \cache_data_reg[14][53]  ( .ip(n4986), .ck(clk), .q(
        \cache_data[14][53] ) );
  dp_1 \cache_data_reg[14][85]  ( .ip(n4954), .ck(clk), .q(
        \cache_data[14][85] ) );
  dp_1 \cache_data_reg[14][117]  ( .ip(n4922), .ck(clk), .q(
        \cache_data[14][117] ) );
  dp_1 \cache_data_reg[15][21]  ( .ip(n4890), .ck(clk), .q(
        \cache_data[15][21] ) );
  dp_1 \cache_data_reg[15][53]  ( .ip(n4858), .ck(clk), .q(
        \cache_data[15][53] ) );
  dp_1 \cache_data_reg[15][85]  ( .ip(n4826), .ck(clk), .q(
        \cache_data[15][85] ) );
  dp_1 \cache_data_reg[15][117]  ( .ip(n4794), .ck(clk), .q(
        \cache_data[15][117] ) );
  dp_1 \iCache_data_wr_reg[22]  ( .ip(n6841), .ck(clk), .q(iCache_data_wr[22])
         );
  dp_1 \cache_data_reg[0][22]  ( .ip(n6809), .ck(clk), .q(\cache_data[0][22] )
         );
  dp_1 \cache_data_reg[0][54]  ( .ip(n6777), .ck(clk), .q(\cache_data[0][54] )
         );
  dp_1 \cache_data_reg[0][86]  ( .ip(n6745), .ck(clk), .q(\cache_data[0][86] )
         );
  dp_1 \cache_data_reg[0][118]  ( .ip(n6713), .ck(clk), .q(
        \cache_data[0][118] ) );
  dp_1 \cache_data_reg[1][22]  ( .ip(n6681), .ck(clk), .q(\cache_data[1][22] )
         );
  dp_1 \cache_data_reg[1][54]  ( .ip(n6649), .ck(clk), .q(\cache_data[1][54] )
         );
  dp_1 \cache_data_reg[1][86]  ( .ip(n6617), .ck(clk), .q(\cache_data[1][86] )
         );
  dp_1 \cache_data_reg[1][118]  ( .ip(n6585), .ck(clk), .q(
        \cache_data[1][118] ) );
  dp_1 \cache_data_reg[2][22]  ( .ip(n6553), .ck(clk), .q(\cache_data[2][22] )
         );
  dp_1 \cache_data_reg[2][54]  ( .ip(n6521), .ck(clk), .q(\cache_data[2][54] )
         );
  dp_1 \cache_data_reg[2][86]  ( .ip(n6489), .ck(clk), .q(\cache_data[2][86] )
         );
  dp_1 \cache_data_reg[2][118]  ( .ip(n6457), .ck(clk), .q(
        \cache_data[2][118] ) );
  dp_1 \cache_data_reg[3][22]  ( .ip(n6425), .ck(clk), .q(\cache_data[3][22] )
         );
  dp_1 \cache_data_reg[3][54]  ( .ip(n6393), .ck(clk), .q(\cache_data[3][54] )
         );
  dp_1 \cache_data_reg[3][86]  ( .ip(n6361), .ck(clk), .q(\cache_data[3][86] )
         );
  dp_1 \cache_data_reg[3][118]  ( .ip(n6329), .ck(clk), .q(
        \cache_data[3][118] ) );
  dp_1 \cache_data_reg[4][22]  ( .ip(n6297), .ck(clk), .q(\cache_data[4][22] )
         );
  dp_1 \cache_data_reg[4][54]  ( .ip(n6265), .ck(clk), .q(\cache_data[4][54] )
         );
  dp_1 \cache_data_reg[4][86]  ( .ip(n6233), .ck(clk), .q(\cache_data[4][86] )
         );
  dp_1 \cache_data_reg[4][118]  ( .ip(n6201), .ck(clk), .q(
        \cache_data[4][118] ) );
  dp_1 \cache_data_reg[5][22]  ( .ip(n6169), .ck(clk), .q(\cache_data[5][22] )
         );
  dp_1 \cache_data_reg[5][54]  ( .ip(n6137), .ck(clk), .q(\cache_data[5][54] )
         );
  dp_1 \cache_data_reg[5][86]  ( .ip(n6105), .ck(clk), .q(\cache_data[5][86] )
         );
  dp_1 \cache_data_reg[5][118]  ( .ip(n6073), .ck(clk), .q(
        \cache_data[5][118] ) );
  dp_1 \cache_data_reg[6][22]  ( .ip(n6041), .ck(clk), .q(\cache_data[6][22] )
         );
  dp_1 \cache_data_reg[6][54]  ( .ip(n6009), .ck(clk), .q(\cache_data[6][54] )
         );
  dp_1 \cache_data_reg[6][86]  ( .ip(n5977), .ck(clk), .q(\cache_data[6][86] )
         );
  dp_1 \cache_data_reg[6][118]  ( .ip(n5945), .ck(clk), .q(
        \cache_data[6][118] ) );
  dp_1 \cache_data_reg[7][22]  ( .ip(n5913), .ck(clk), .q(\cache_data[7][22] )
         );
  dp_1 \cache_data_reg[7][54]  ( .ip(n5881), .ck(clk), .q(\cache_data[7][54] )
         );
  dp_1 \cache_data_reg[7][86]  ( .ip(n5849), .ck(clk), .q(\cache_data[7][86] )
         );
  dp_1 \cache_data_reg[7][118]  ( .ip(n5817), .ck(clk), .q(
        \cache_data[7][118] ) );
  dp_1 \cache_data_reg[8][22]  ( .ip(n5785), .ck(clk), .q(\cache_data[8][22] )
         );
  dp_1 \cache_data_reg[8][54]  ( .ip(n5753), .ck(clk), .q(\cache_data[8][54] )
         );
  dp_1 \cache_data_reg[8][86]  ( .ip(n5721), .ck(clk), .q(\cache_data[8][86] )
         );
  dp_1 \cache_data_reg[8][118]  ( .ip(n5689), .ck(clk), .q(
        \cache_data[8][118] ) );
  dp_1 \cache_data_reg[9][22]  ( .ip(n5657), .ck(clk), .q(\cache_data[9][22] )
         );
  dp_1 \cache_data_reg[9][54]  ( .ip(n5625), .ck(clk), .q(\cache_data[9][54] )
         );
  dp_1 \cache_data_reg[9][86]  ( .ip(n5593), .ck(clk), .q(\cache_data[9][86] )
         );
  dp_1 \cache_data_reg[9][118]  ( .ip(n5561), .ck(clk), .q(
        \cache_data[9][118] ) );
  dp_1 \cache_data_reg[10][22]  ( .ip(n5529), .ck(clk), .q(
        \cache_data[10][22] ) );
  dp_1 \cache_data_reg[10][54]  ( .ip(n5497), .ck(clk), .q(
        \cache_data[10][54] ) );
  dp_1 \cache_data_reg[10][86]  ( .ip(n5465), .ck(clk), .q(
        \cache_data[10][86] ) );
  dp_1 \cache_data_reg[10][118]  ( .ip(n5433), .ck(clk), .q(
        \cache_data[10][118] ) );
  dp_1 \cache_data_reg[11][22]  ( .ip(n5401), .ck(clk), .q(
        \cache_data[11][22] ) );
  dp_1 \cache_data_reg[11][54]  ( .ip(n5369), .ck(clk), .q(
        \cache_data[11][54] ) );
  dp_1 \cache_data_reg[11][86]  ( .ip(n5337), .ck(clk), .q(
        \cache_data[11][86] ) );
  dp_1 \cache_data_reg[11][118]  ( .ip(n5305), .ck(clk), .q(
        \cache_data[11][118] ) );
  dp_1 \cache_data_reg[12][22]  ( .ip(n5273), .ck(clk), .q(
        \cache_data[12][22] ) );
  dp_1 \cache_data_reg[12][54]  ( .ip(n5241), .ck(clk), .q(
        \cache_data[12][54] ) );
  dp_1 \cache_data_reg[12][86]  ( .ip(n5209), .ck(clk), .q(
        \cache_data[12][86] ) );
  dp_1 \cache_data_reg[12][118]  ( .ip(n5177), .ck(clk), .q(
        \cache_data[12][118] ) );
  dp_1 \cache_data_reg[13][22]  ( .ip(n5145), .ck(clk), .q(
        \cache_data[13][22] ) );
  dp_1 \cache_data_reg[13][54]  ( .ip(n5113), .ck(clk), .q(
        \cache_data[13][54] ) );
  dp_1 \cache_data_reg[13][86]  ( .ip(n5081), .ck(clk), .q(
        \cache_data[13][86] ) );
  dp_1 \cache_data_reg[13][118]  ( .ip(n5049), .ck(clk), .q(
        \cache_data[13][118] ) );
  dp_1 \cache_data_reg[14][22]  ( .ip(n5017), .ck(clk), .q(
        \cache_data[14][22] ) );
  dp_1 \cache_data_reg[14][54]  ( .ip(n4985), .ck(clk), .q(
        \cache_data[14][54] ) );
  dp_1 \cache_data_reg[14][86]  ( .ip(n4953), .ck(clk), .q(
        \cache_data[14][86] ) );
  dp_1 \cache_data_reg[14][118]  ( .ip(n4921), .ck(clk), .q(
        \cache_data[14][118] ) );
  dp_1 \cache_data_reg[15][22]  ( .ip(n4889), .ck(clk), .q(
        \cache_data[15][22] ) );
  dp_1 \cache_data_reg[15][54]  ( .ip(n4857), .ck(clk), .q(
        \cache_data[15][54] ) );
  dp_1 \cache_data_reg[15][86]  ( .ip(n4825), .ck(clk), .q(
        \cache_data[15][86] ) );
  dp_1 \cache_data_reg[15][118]  ( .ip(n4793), .ck(clk), .q(
        \cache_data[15][118] ) );
  dp_1 \iCache_data_wr_reg[23]  ( .ip(n6840), .ck(clk), .q(iCache_data_wr[23])
         );
  dp_1 \cache_data_reg[0][23]  ( .ip(n6808), .ck(clk), .q(\cache_data[0][23] )
         );
  dp_1 \cache_data_reg[0][55]  ( .ip(n6776), .ck(clk), .q(\cache_data[0][55] )
         );
  dp_1 \cache_data_reg[0][87]  ( .ip(n6744), .ck(clk), .q(\cache_data[0][87] )
         );
  dp_1 \cache_data_reg[0][119]  ( .ip(n6712), .ck(clk), .q(
        \cache_data[0][119] ) );
  dp_1 \cache_data_reg[1][23]  ( .ip(n6680), .ck(clk), .q(\cache_data[1][23] )
         );
  dp_1 \cache_data_reg[1][55]  ( .ip(n6648), .ck(clk), .q(\cache_data[1][55] )
         );
  dp_1 \cache_data_reg[1][87]  ( .ip(n6616), .ck(clk), .q(\cache_data[1][87] )
         );
  dp_1 \cache_data_reg[1][119]  ( .ip(n6584), .ck(clk), .q(
        \cache_data[1][119] ) );
  dp_1 \cache_data_reg[2][23]  ( .ip(n6552), .ck(clk), .q(\cache_data[2][23] )
         );
  dp_1 \cache_data_reg[2][55]  ( .ip(n6520), .ck(clk), .q(\cache_data[2][55] )
         );
  dp_1 \cache_data_reg[2][87]  ( .ip(n6488), .ck(clk), .q(\cache_data[2][87] )
         );
  dp_1 \cache_data_reg[2][119]  ( .ip(n6456), .ck(clk), .q(
        \cache_data[2][119] ) );
  dp_1 \cache_data_reg[3][23]  ( .ip(n6424), .ck(clk), .q(\cache_data[3][23] )
         );
  dp_1 \cache_data_reg[3][55]  ( .ip(n6392), .ck(clk), .q(\cache_data[3][55] )
         );
  dp_1 \cache_data_reg[3][87]  ( .ip(n6360), .ck(clk), .q(\cache_data[3][87] )
         );
  dp_1 \cache_data_reg[3][119]  ( .ip(n6328), .ck(clk), .q(
        \cache_data[3][119] ) );
  dp_1 \cache_data_reg[4][23]  ( .ip(n6296), .ck(clk), .q(\cache_data[4][23] )
         );
  dp_1 \cache_data_reg[4][55]  ( .ip(n6264), .ck(clk), .q(\cache_data[4][55] )
         );
  dp_1 \cache_data_reg[4][87]  ( .ip(n6232), .ck(clk), .q(\cache_data[4][87] )
         );
  dp_1 \cache_data_reg[4][119]  ( .ip(n6200), .ck(clk), .q(
        \cache_data[4][119] ) );
  dp_1 \cache_data_reg[5][23]  ( .ip(n6168), .ck(clk), .q(\cache_data[5][23] )
         );
  dp_1 \cache_data_reg[5][55]  ( .ip(n6136), .ck(clk), .q(\cache_data[5][55] )
         );
  dp_1 \cache_data_reg[5][87]  ( .ip(n6104), .ck(clk), .q(\cache_data[5][87] )
         );
  dp_1 \cache_data_reg[5][119]  ( .ip(n6072), .ck(clk), .q(
        \cache_data[5][119] ) );
  dp_1 \cache_data_reg[6][23]  ( .ip(n6040), .ck(clk), .q(\cache_data[6][23] )
         );
  dp_1 \cache_data_reg[6][55]  ( .ip(n6008), .ck(clk), .q(\cache_data[6][55] )
         );
  dp_1 \cache_data_reg[6][87]  ( .ip(n5976), .ck(clk), .q(\cache_data[6][87] )
         );
  dp_1 \cache_data_reg[6][119]  ( .ip(n5944), .ck(clk), .q(
        \cache_data[6][119] ) );
  dp_1 \cache_data_reg[7][23]  ( .ip(n5912), .ck(clk), .q(\cache_data[7][23] )
         );
  dp_1 \cache_data_reg[7][55]  ( .ip(n5880), .ck(clk), .q(\cache_data[7][55] )
         );
  dp_1 \cache_data_reg[7][87]  ( .ip(n5848), .ck(clk), .q(\cache_data[7][87] )
         );
  dp_1 \cache_data_reg[7][119]  ( .ip(n5816), .ck(clk), .q(
        \cache_data[7][119] ) );
  dp_1 \cache_data_reg[8][23]  ( .ip(n5784), .ck(clk), .q(\cache_data[8][23] )
         );
  dp_1 \cache_data_reg[8][55]  ( .ip(n5752), .ck(clk), .q(\cache_data[8][55] )
         );
  dp_1 \cache_data_reg[8][87]  ( .ip(n5720), .ck(clk), .q(\cache_data[8][87] )
         );
  dp_1 \cache_data_reg[8][119]  ( .ip(n5688), .ck(clk), .q(
        \cache_data[8][119] ) );
  dp_1 \cache_data_reg[9][23]  ( .ip(n5656), .ck(clk), .q(\cache_data[9][23] )
         );
  dp_1 \cache_data_reg[9][55]  ( .ip(n5624), .ck(clk), .q(\cache_data[9][55] )
         );
  dp_1 \cache_data_reg[9][87]  ( .ip(n5592), .ck(clk), .q(\cache_data[9][87] )
         );
  dp_1 \cache_data_reg[9][119]  ( .ip(n5560), .ck(clk), .q(
        \cache_data[9][119] ) );
  dp_1 \cache_data_reg[10][23]  ( .ip(n5528), .ck(clk), .q(
        \cache_data[10][23] ) );
  dp_1 \cache_data_reg[10][55]  ( .ip(n5496), .ck(clk), .q(
        \cache_data[10][55] ) );
  dp_1 \cache_data_reg[10][87]  ( .ip(n5464), .ck(clk), .q(
        \cache_data[10][87] ) );
  dp_1 \cache_data_reg[10][119]  ( .ip(n5432), .ck(clk), .q(
        \cache_data[10][119] ) );
  dp_1 \cache_data_reg[11][23]  ( .ip(n5400), .ck(clk), .q(
        \cache_data[11][23] ) );
  dp_1 \cache_data_reg[11][55]  ( .ip(n5368), .ck(clk), .q(
        \cache_data[11][55] ) );
  dp_1 \cache_data_reg[11][87]  ( .ip(n5336), .ck(clk), .q(
        \cache_data[11][87] ) );
  dp_1 \cache_data_reg[11][119]  ( .ip(n5304), .ck(clk), .q(
        \cache_data[11][119] ) );
  dp_1 \cache_data_reg[12][23]  ( .ip(n5272), .ck(clk), .q(
        \cache_data[12][23] ) );
  dp_1 \cache_data_reg[12][55]  ( .ip(n5240), .ck(clk), .q(
        \cache_data[12][55] ) );
  dp_1 \cache_data_reg[12][87]  ( .ip(n5208), .ck(clk), .q(
        \cache_data[12][87] ) );
  dp_1 \cache_data_reg[12][119]  ( .ip(n5176), .ck(clk), .q(
        \cache_data[12][119] ) );
  dp_1 \cache_data_reg[13][23]  ( .ip(n5144), .ck(clk), .q(
        \cache_data[13][23] ) );
  dp_1 \cache_data_reg[13][55]  ( .ip(n5112), .ck(clk), .q(
        \cache_data[13][55] ) );
  dp_1 \cache_data_reg[13][87]  ( .ip(n5080), .ck(clk), .q(
        \cache_data[13][87] ) );
  dp_1 \cache_data_reg[13][119]  ( .ip(n5048), .ck(clk), .q(
        \cache_data[13][119] ) );
  dp_1 \cache_data_reg[14][23]  ( .ip(n5016), .ck(clk), .q(
        \cache_data[14][23] ) );
  dp_1 \cache_data_reg[14][55]  ( .ip(n4984), .ck(clk), .q(
        \cache_data[14][55] ) );
  dp_1 \cache_data_reg[14][87]  ( .ip(n4952), .ck(clk), .q(
        \cache_data[14][87] ) );
  dp_1 \cache_data_reg[14][119]  ( .ip(n4920), .ck(clk), .q(
        \cache_data[14][119] ) );
  dp_1 \cache_data_reg[15][23]  ( .ip(n4888), .ck(clk), .q(
        \cache_data[15][23] ) );
  dp_1 \cache_data_reg[15][55]  ( .ip(n4856), .ck(clk), .q(
        \cache_data[15][55] ) );
  dp_1 \cache_data_reg[15][87]  ( .ip(n4824), .ck(clk), .q(
        \cache_data[15][87] ) );
  dp_1 \cache_data_reg[15][119]  ( .ip(n4792), .ck(clk), .q(
        \cache_data[15][119] ) );
  dp_1 \iCache_data_wr_reg[24]  ( .ip(n6839), .ck(clk), .q(iCache_data_wr[24])
         );
  dp_1 \cache_data_reg[0][24]  ( .ip(n6807), .ck(clk), .q(\cache_data[0][24] )
         );
  dp_1 \cache_data_reg[0][56]  ( .ip(n6775), .ck(clk), .q(\cache_data[0][56] )
         );
  dp_1 \cache_data_reg[0][88]  ( .ip(n6743), .ck(clk), .q(\cache_data[0][88] )
         );
  dp_1 \cache_data_reg[0][120]  ( .ip(n6711), .ck(clk), .q(
        \cache_data[0][120] ) );
  dp_1 \cache_data_reg[1][24]  ( .ip(n6679), .ck(clk), .q(\cache_data[1][24] )
         );
  dp_1 \cache_data_reg[1][56]  ( .ip(n6647), .ck(clk), .q(\cache_data[1][56] )
         );
  dp_1 \cache_data_reg[1][88]  ( .ip(n6615), .ck(clk), .q(\cache_data[1][88] )
         );
  dp_1 \cache_data_reg[1][120]  ( .ip(n6583), .ck(clk), .q(
        \cache_data[1][120] ) );
  dp_1 \cache_data_reg[2][24]  ( .ip(n6551), .ck(clk), .q(\cache_data[2][24] )
         );
  dp_1 \cache_data_reg[2][56]  ( .ip(n6519), .ck(clk), .q(\cache_data[2][56] )
         );
  dp_1 \cache_data_reg[2][88]  ( .ip(n6487), .ck(clk), .q(\cache_data[2][88] )
         );
  dp_1 \cache_data_reg[2][120]  ( .ip(n6455), .ck(clk), .q(
        \cache_data[2][120] ) );
  dp_1 \cache_data_reg[3][24]  ( .ip(n6423), .ck(clk), .q(\cache_data[3][24] )
         );
  dp_1 \cache_data_reg[3][56]  ( .ip(n6391), .ck(clk), .q(\cache_data[3][56] )
         );
  dp_1 \cache_data_reg[3][88]  ( .ip(n6359), .ck(clk), .q(\cache_data[3][88] )
         );
  dp_1 \cache_data_reg[3][120]  ( .ip(n6327), .ck(clk), .q(
        \cache_data[3][120] ) );
  dp_1 \cache_data_reg[4][24]  ( .ip(n6295), .ck(clk), .q(\cache_data[4][24] )
         );
  dp_1 \cache_data_reg[4][56]  ( .ip(n6263), .ck(clk), .q(\cache_data[4][56] )
         );
  dp_1 \cache_data_reg[4][88]  ( .ip(n6231), .ck(clk), .q(\cache_data[4][88] )
         );
  dp_1 \cache_data_reg[4][120]  ( .ip(n6199), .ck(clk), .q(
        \cache_data[4][120] ) );
  dp_1 \cache_data_reg[5][24]  ( .ip(n6167), .ck(clk), .q(\cache_data[5][24] )
         );
  dp_1 \cache_data_reg[5][56]  ( .ip(n6135), .ck(clk), .q(\cache_data[5][56] )
         );
  dp_1 \cache_data_reg[5][88]  ( .ip(n6103), .ck(clk), .q(\cache_data[5][88] )
         );
  dp_1 \cache_data_reg[5][120]  ( .ip(n6071), .ck(clk), .q(
        \cache_data[5][120] ) );
  dp_1 \cache_data_reg[6][24]  ( .ip(n6039), .ck(clk), .q(\cache_data[6][24] )
         );
  dp_1 \cache_data_reg[6][56]  ( .ip(n6007), .ck(clk), .q(\cache_data[6][56] )
         );
  dp_1 \cache_data_reg[6][88]  ( .ip(n5975), .ck(clk), .q(\cache_data[6][88] )
         );
  dp_1 \cache_data_reg[6][120]  ( .ip(n5943), .ck(clk), .q(
        \cache_data[6][120] ) );
  dp_1 \cache_data_reg[7][24]  ( .ip(n5911), .ck(clk), .q(\cache_data[7][24] )
         );
  dp_1 \cache_data_reg[7][56]  ( .ip(n5879), .ck(clk), .q(\cache_data[7][56] )
         );
  dp_1 \cache_data_reg[7][88]  ( .ip(n5847), .ck(clk), .q(\cache_data[7][88] )
         );
  dp_1 \cache_data_reg[7][120]  ( .ip(n5815), .ck(clk), .q(
        \cache_data[7][120] ) );
  dp_1 \cache_data_reg[8][24]  ( .ip(n5783), .ck(clk), .q(\cache_data[8][24] )
         );
  dp_1 \cache_data_reg[8][56]  ( .ip(n5751), .ck(clk), .q(\cache_data[8][56] )
         );
  dp_1 \cache_data_reg[8][88]  ( .ip(n5719), .ck(clk), .q(\cache_data[8][88] )
         );
  dp_1 \cache_data_reg[8][120]  ( .ip(n5687), .ck(clk), .q(
        \cache_data[8][120] ) );
  dp_1 \cache_data_reg[9][24]  ( .ip(n5655), .ck(clk), .q(\cache_data[9][24] )
         );
  dp_1 \cache_data_reg[9][56]  ( .ip(n5623), .ck(clk), .q(\cache_data[9][56] )
         );
  dp_1 \cache_data_reg[9][88]  ( .ip(n5591), .ck(clk), .q(\cache_data[9][88] )
         );
  dp_1 \cache_data_reg[9][120]  ( .ip(n5559), .ck(clk), .q(
        \cache_data[9][120] ) );
  dp_1 \cache_data_reg[10][24]  ( .ip(n5527), .ck(clk), .q(
        \cache_data[10][24] ) );
  dp_1 \cache_data_reg[10][56]  ( .ip(n5495), .ck(clk), .q(
        \cache_data[10][56] ) );
  dp_1 \cache_data_reg[10][88]  ( .ip(n5463), .ck(clk), .q(
        \cache_data[10][88] ) );
  dp_1 \cache_data_reg[10][120]  ( .ip(n5431), .ck(clk), .q(
        \cache_data[10][120] ) );
  dp_1 \cache_data_reg[11][24]  ( .ip(n5399), .ck(clk), .q(
        \cache_data[11][24] ) );
  dp_1 \cache_data_reg[11][56]  ( .ip(n5367), .ck(clk), .q(
        \cache_data[11][56] ) );
  dp_1 \cache_data_reg[11][88]  ( .ip(n5335), .ck(clk), .q(
        \cache_data[11][88] ) );
  dp_1 \cache_data_reg[11][120]  ( .ip(n5303), .ck(clk), .q(
        \cache_data[11][120] ) );
  dp_1 \cache_data_reg[12][24]  ( .ip(n5271), .ck(clk), .q(
        \cache_data[12][24] ) );
  dp_1 \cache_data_reg[12][56]  ( .ip(n5239), .ck(clk), .q(
        \cache_data[12][56] ) );
  dp_1 \cache_data_reg[12][88]  ( .ip(n5207), .ck(clk), .q(
        \cache_data[12][88] ) );
  dp_1 \cache_data_reg[12][120]  ( .ip(n5175), .ck(clk), .q(
        \cache_data[12][120] ) );
  dp_1 \cache_data_reg[13][24]  ( .ip(n5143), .ck(clk), .q(
        \cache_data[13][24] ) );
  dp_1 \cache_data_reg[13][56]  ( .ip(n5111), .ck(clk), .q(
        \cache_data[13][56] ) );
  dp_1 \cache_data_reg[13][88]  ( .ip(n5079), .ck(clk), .q(
        \cache_data[13][88] ) );
  dp_1 \cache_data_reg[13][120]  ( .ip(n5047), .ck(clk), .q(
        \cache_data[13][120] ) );
  dp_1 \cache_data_reg[14][24]  ( .ip(n5015), .ck(clk), .q(
        \cache_data[14][24] ) );
  dp_1 \cache_data_reg[14][56]  ( .ip(n4983), .ck(clk), .q(
        \cache_data[14][56] ) );
  dp_1 \cache_data_reg[14][88]  ( .ip(n4951), .ck(clk), .q(
        \cache_data[14][88] ) );
  dp_1 \cache_data_reg[14][120]  ( .ip(n4919), .ck(clk), .q(
        \cache_data[14][120] ) );
  dp_1 \cache_data_reg[15][24]  ( .ip(n4887), .ck(clk), .q(
        \cache_data[15][24] ) );
  dp_1 \cache_data_reg[15][56]  ( .ip(n4855), .ck(clk), .q(
        \cache_data[15][56] ) );
  dp_1 \cache_data_reg[15][88]  ( .ip(n4823), .ck(clk), .q(
        \cache_data[15][88] ) );
  dp_1 \cache_data_reg[15][120]  ( .ip(n4791), .ck(clk), .q(
        \cache_data[15][120] ) );
  dp_1 \iCache_data_wr_reg[25]  ( .ip(n6838), .ck(clk), .q(iCache_data_wr[25])
         );
  dp_1 \cache_data_reg[0][25]  ( .ip(n6806), .ck(clk), .q(\cache_data[0][25] )
         );
  dp_1 \cache_data_reg[0][57]  ( .ip(n6774), .ck(clk), .q(\cache_data[0][57] )
         );
  dp_1 \cache_data_reg[0][89]  ( .ip(n6742), .ck(clk), .q(\cache_data[0][89] )
         );
  dp_1 \cache_data_reg[0][121]  ( .ip(n6710), .ck(clk), .q(
        \cache_data[0][121] ) );
  dp_1 \cache_data_reg[1][25]  ( .ip(n6678), .ck(clk), .q(\cache_data[1][25] )
         );
  dp_1 \cache_data_reg[1][57]  ( .ip(n6646), .ck(clk), .q(\cache_data[1][57] )
         );
  dp_1 \cache_data_reg[1][89]  ( .ip(n6614), .ck(clk), .q(\cache_data[1][89] )
         );
  dp_1 \cache_data_reg[1][121]  ( .ip(n6582), .ck(clk), .q(
        \cache_data[1][121] ) );
  dp_1 \cache_data_reg[2][25]  ( .ip(n6550), .ck(clk), .q(\cache_data[2][25] )
         );
  dp_1 \cache_data_reg[2][57]  ( .ip(n6518), .ck(clk), .q(\cache_data[2][57] )
         );
  dp_1 \cache_data_reg[2][89]  ( .ip(n6486), .ck(clk), .q(\cache_data[2][89] )
         );
  dp_1 \cache_data_reg[2][121]  ( .ip(n6454), .ck(clk), .q(
        \cache_data[2][121] ) );
  dp_1 \cache_data_reg[3][25]  ( .ip(n6422), .ck(clk), .q(\cache_data[3][25] )
         );
  dp_1 \cache_data_reg[3][57]  ( .ip(n6390), .ck(clk), .q(\cache_data[3][57] )
         );
  dp_1 \cache_data_reg[3][89]  ( .ip(n6358), .ck(clk), .q(\cache_data[3][89] )
         );
  dp_1 \cache_data_reg[3][121]  ( .ip(n6326), .ck(clk), .q(
        \cache_data[3][121] ) );
  dp_1 \cache_data_reg[4][25]  ( .ip(n6294), .ck(clk), .q(\cache_data[4][25] )
         );
  dp_1 \cache_data_reg[4][57]  ( .ip(n6262), .ck(clk), .q(\cache_data[4][57] )
         );
  dp_1 \cache_data_reg[4][89]  ( .ip(n6230), .ck(clk), .q(\cache_data[4][89] )
         );
  dp_1 \cache_data_reg[4][121]  ( .ip(n6198), .ck(clk), .q(
        \cache_data[4][121] ) );
  dp_1 \cache_data_reg[5][25]  ( .ip(n6166), .ck(clk), .q(\cache_data[5][25] )
         );
  dp_1 \cache_data_reg[5][57]  ( .ip(n6134), .ck(clk), .q(\cache_data[5][57] )
         );
  dp_1 \cache_data_reg[5][89]  ( .ip(n6102), .ck(clk), .q(\cache_data[5][89] )
         );
  dp_1 \cache_data_reg[5][121]  ( .ip(n6070), .ck(clk), .q(
        \cache_data[5][121] ) );
  dp_1 \cache_data_reg[6][25]  ( .ip(n6038), .ck(clk), .q(\cache_data[6][25] )
         );
  dp_1 \cache_data_reg[6][57]  ( .ip(n6006), .ck(clk), .q(\cache_data[6][57] )
         );
  dp_1 \cache_data_reg[6][89]  ( .ip(n5974), .ck(clk), .q(\cache_data[6][89] )
         );
  dp_1 \cache_data_reg[6][121]  ( .ip(n5942), .ck(clk), .q(
        \cache_data[6][121] ) );
  dp_1 \cache_data_reg[7][25]  ( .ip(n5910), .ck(clk), .q(\cache_data[7][25] )
         );
  dp_1 \cache_data_reg[7][57]  ( .ip(n5878), .ck(clk), .q(\cache_data[7][57] )
         );
  dp_1 \cache_data_reg[7][89]  ( .ip(n5846), .ck(clk), .q(\cache_data[7][89] )
         );
  dp_1 \cache_data_reg[7][121]  ( .ip(n5814), .ck(clk), .q(
        \cache_data[7][121] ) );
  dp_1 \cache_data_reg[8][25]  ( .ip(n5782), .ck(clk), .q(\cache_data[8][25] )
         );
  dp_1 \cache_data_reg[8][57]  ( .ip(n5750), .ck(clk), .q(\cache_data[8][57] )
         );
  dp_1 \cache_data_reg[8][89]  ( .ip(n5718), .ck(clk), .q(\cache_data[8][89] )
         );
  dp_1 \cache_data_reg[8][121]  ( .ip(n5686), .ck(clk), .q(
        \cache_data[8][121] ) );
  dp_1 \cache_data_reg[9][25]  ( .ip(n5654), .ck(clk), .q(\cache_data[9][25] )
         );
  dp_1 \cache_data_reg[9][57]  ( .ip(n5622), .ck(clk), .q(\cache_data[9][57] )
         );
  dp_1 \cache_data_reg[9][89]  ( .ip(n5590), .ck(clk), .q(\cache_data[9][89] )
         );
  dp_1 \cache_data_reg[9][121]  ( .ip(n5558), .ck(clk), .q(
        \cache_data[9][121] ) );
  dp_1 \cache_data_reg[10][25]  ( .ip(n5526), .ck(clk), .q(
        \cache_data[10][25] ) );
  dp_1 \cache_data_reg[10][57]  ( .ip(n5494), .ck(clk), .q(
        \cache_data[10][57] ) );
  dp_1 \cache_data_reg[10][89]  ( .ip(n5462), .ck(clk), .q(
        \cache_data[10][89] ) );
  dp_1 \cache_data_reg[10][121]  ( .ip(n5430), .ck(clk), .q(
        \cache_data[10][121] ) );
  dp_1 \cache_data_reg[11][25]  ( .ip(n5398), .ck(clk), .q(
        \cache_data[11][25] ) );
  dp_1 \cache_data_reg[11][57]  ( .ip(n5366), .ck(clk), .q(
        \cache_data[11][57] ) );
  dp_1 \cache_data_reg[11][89]  ( .ip(n5334), .ck(clk), .q(
        \cache_data[11][89] ) );
  dp_1 \cache_data_reg[11][121]  ( .ip(n5302), .ck(clk), .q(
        \cache_data[11][121] ) );
  dp_1 \cache_data_reg[12][25]  ( .ip(n5270), .ck(clk), .q(
        \cache_data[12][25] ) );
  dp_1 \cache_data_reg[12][57]  ( .ip(n5238), .ck(clk), .q(
        \cache_data[12][57] ) );
  dp_1 \cache_data_reg[12][89]  ( .ip(n5206), .ck(clk), .q(
        \cache_data[12][89] ) );
  dp_1 \cache_data_reg[12][121]  ( .ip(n5174), .ck(clk), .q(
        \cache_data[12][121] ) );
  dp_1 \cache_data_reg[13][25]  ( .ip(n5142), .ck(clk), .q(
        \cache_data[13][25] ) );
  dp_1 \cache_data_reg[13][57]  ( .ip(n5110), .ck(clk), .q(
        \cache_data[13][57] ) );
  dp_1 \cache_data_reg[13][89]  ( .ip(n5078), .ck(clk), .q(
        \cache_data[13][89] ) );
  dp_1 \cache_data_reg[13][121]  ( .ip(n5046), .ck(clk), .q(
        \cache_data[13][121] ) );
  dp_1 \cache_data_reg[14][25]  ( .ip(n5014), .ck(clk), .q(
        \cache_data[14][25] ) );
  dp_1 \cache_data_reg[14][57]  ( .ip(n4982), .ck(clk), .q(
        \cache_data[14][57] ) );
  dp_1 \cache_data_reg[14][89]  ( .ip(n4950), .ck(clk), .q(
        \cache_data[14][89] ) );
  dp_1 \cache_data_reg[14][121]  ( .ip(n4918), .ck(clk), .q(
        \cache_data[14][121] ) );
  dp_1 \cache_data_reg[15][25]  ( .ip(n4886), .ck(clk), .q(
        \cache_data[15][25] ) );
  dp_1 \cache_data_reg[15][57]  ( .ip(n4854), .ck(clk), .q(
        \cache_data[15][57] ) );
  dp_1 \cache_data_reg[15][89]  ( .ip(n4822), .ck(clk), .q(
        \cache_data[15][89] ) );
  dp_1 \cache_data_reg[15][121]  ( .ip(n4790), .ck(clk), .q(
        \cache_data[15][121] ) );
  dp_1 \iCache_data_wr_reg[26]  ( .ip(n6837), .ck(clk), .q(iCache_data_wr[26])
         );
  dp_1 \cache_data_reg[0][26]  ( .ip(n6805), .ck(clk), .q(\cache_data[0][26] )
         );
  dp_1 \cache_data_reg[0][58]  ( .ip(n6773), .ck(clk), .q(\cache_data[0][58] )
         );
  dp_1 \cache_data_reg[0][90]  ( .ip(n6741), .ck(clk), .q(\cache_data[0][90] )
         );
  dp_1 \cache_data_reg[0][122]  ( .ip(n6709), .ck(clk), .q(
        \cache_data[0][122] ) );
  dp_1 \cache_data_reg[1][26]  ( .ip(n6677), .ck(clk), .q(\cache_data[1][26] )
         );
  dp_1 \cache_data_reg[1][58]  ( .ip(n6645), .ck(clk), .q(\cache_data[1][58] )
         );
  dp_1 \cache_data_reg[1][90]  ( .ip(n6613), .ck(clk), .q(\cache_data[1][90] )
         );
  dp_1 \cache_data_reg[1][122]  ( .ip(n6581), .ck(clk), .q(
        \cache_data[1][122] ) );
  dp_1 \cache_data_reg[2][26]  ( .ip(n6549), .ck(clk), .q(\cache_data[2][26] )
         );
  dp_1 \cache_data_reg[2][58]  ( .ip(n6517), .ck(clk), .q(\cache_data[2][58] )
         );
  dp_1 \cache_data_reg[2][90]  ( .ip(n6485), .ck(clk), .q(\cache_data[2][90] )
         );
  dp_1 \cache_data_reg[2][122]  ( .ip(n6453), .ck(clk), .q(
        \cache_data[2][122] ) );
  dp_1 \cache_data_reg[3][26]  ( .ip(n6421), .ck(clk), .q(\cache_data[3][26] )
         );
  dp_1 \cache_data_reg[3][58]  ( .ip(n6389), .ck(clk), .q(\cache_data[3][58] )
         );
  dp_1 \cache_data_reg[3][90]  ( .ip(n6357), .ck(clk), .q(\cache_data[3][90] )
         );
  dp_1 \cache_data_reg[3][122]  ( .ip(n6325), .ck(clk), .q(
        \cache_data[3][122] ) );
  dp_1 \cache_data_reg[4][26]  ( .ip(n6293), .ck(clk), .q(\cache_data[4][26] )
         );
  dp_1 \cache_data_reg[4][58]  ( .ip(n6261), .ck(clk), .q(\cache_data[4][58] )
         );
  dp_1 \cache_data_reg[4][90]  ( .ip(n6229), .ck(clk), .q(\cache_data[4][90] )
         );
  dp_1 \cache_data_reg[4][122]  ( .ip(n6197), .ck(clk), .q(
        \cache_data[4][122] ) );
  dp_1 \cache_data_reg[5][26]  ( .ip(n6165), .ck(clk), .q(\cache_data[5][26] )
         );
  dp_1 \cache_data_reg[5][58]  ( .ip(n6133), .ck(clk), .q(\cache_data[5][58] )
         );
  dp_1 \cache_data_reg[5][90]  ( .ip(n6101), .ck(clk), .q(\cache_data[5][90] )
         );
  dp_1 \cache_data_reg[5][122]  ( .ip(n6069), .ck(clk), .q(
        \cache_data[5][122] ) );
  dp_1 \cache_data_reg[6][26]  ( .ip(n6037), .ck(clk), .q(\cache_data[6][26] )
         );
  dp_1 \cache_data_reg[6][58]  ( .ip(n6005), .ck(clk), .q(\cache_data[6][58] )
         );
  dp_1 \cache_data_reg[6][90]  ( .ip(n5973), .ck(clk), .q(\cache_data[6][90] )
         );
  dp_1 \cache_data_reg[6][122]  ( .ip(n5941), .ck(clk), .q(
        \cache_data[6][122] ) );
  dp_1 \cache_data_reg[7][26]  ( .ip(n5909), .ck(clk), .q(\cache_data[7][26] )
         );
  dp_1 \cache_data_reg[7][58]  ( .ip(n5877), .ck(clk), .q(\cache_data[7][58] )
         );
  dp_1 \cache_data_reg[7][90]  ( .ip(n5845), .ck(clk), .q(\cache_data[7][90] )
         );
  dp_1 \cache_data_reg[7][122]  ( .ip(n5813), .ck(clk), .q(
        \cache_data[7][122] ) );
  dp_1 \cache_data_reg[8][26]  ( .ip(n5781), .ck(clk), .q(\cache_data[8][26] )
         );
  dp_1 \cache_data_reg[8][58]  ( .ip(n5749), .ck(clk), .q(\cache_data[8][58] )
         );
  dp_1 \cache_data_reg[8][90]  ( .ip(n5717), .ck(clk), .q(\cache_data[8][90] )
         );
  dp_1 \cache_data_reg[8][122]  ( .ip(n5685), .ck(clk), .q(
        \cache_data[8][122] ) );
  dp_1 \cache_data_reg[9][26]  ( .ip(n5653), .ck(clk), .q(\cache_data[9][26] )
         );
  dp_1 \cache_data_reg[9][58]  ( .ip(n5621), .ck(clk), .q(\cache_data[9][58] )
         );
  dp_1 \cache_data_reg[9][90]  ( .ip(n5589), .ck(clk), .q(\cache_data[9][90] )
         );
  dp_1 \cache_data_reg[9][122]  ( .ip(n5557), .ck(clk), .q(
        \cache_data[9][122] ) );
  dp_1 \cache_data_reg[10][26]  ( .ip(n5525), .ck(clk), .q(
        \cache_data[10][26] ) );
  dp_1 \cache_data_reg[10][58]  ( .ip(n5493), .ck(clk), .q(
        \cache_data[10][58] ) );
  dp_1 \cache_data_reg[10][90]  ( .ip(n5461), .ck(clk), .q(
        \cache_data[10][90] ) );
  dp_1 \cache_data_reg[10][122]  ( .ip(n5429), .ck(clk), .q(
        \cache_data[10][122] ) );
  dp_1 \cache_data_reg[11][26]  ( .ip(n5397), .ck(clk), .q(
        \cache_data[11][26] ) );
  dp_1 \cache_data_reg[11][58]  ( .ip(n5365), .ck(clk), .q(
        \cache_data[11][58] ) );
  dp_1 \cache_data_reg[11][90]  ( .ip(n5333), .ck(clk), .q(
        \cache_data[11][90] ) );
  dp_1 \cache_data_reg[11][122]  ( .ip(n5301), .ck(clk), .q(
        \cache_data[11][122] ) );
  dp_1 \cache_data_reg[12][26]  ( .ip(n5269), .ck(clk), .q(
        \cache_data[12][26] ) );
  dp_1 \cache_data_reg[12][58]  ( .ip(n5237), .ck(clk), .q(
        \cache_data[12][58] ) );
  dp_1 \cache_data_reg[12][90]  ( .ip(n5205), .ck(clk), .q(
        \cache_data[12][90] ) );
  dp_1 \cache_data_reg[12][122]  ( .ip(n5173), .ck(clk), .q(
        \cache_data[12][122] ) );
  dp_1 \cache_data_reg[13][26]  ( .ip(n5141), .ck(clk), .q(
        \cache_data[13][26] ) );
  dp_1 \cache_data_reg[13][58]  ( .ip(n5109), .ck(clk), .q(
        \cache_data[13][58] ) );
  dp_1 \cache_data_reg[13][90]  ( .ip(n5077), .ck(clk), .q(
        \cache_data[13][90] ) );
  dp_1 \cache_data_reg[13][122]  ( .ip(n5045), .ck(clk), .q(
        \cache_data[13][122] ) );
  dp_1 \cache_data_reg[14][26]  ( .ip(n5013), .ck(clk), .q(
        \cache_data[14][26] ) );
  dp_1 \cache_data_reg[14][58]  ( .ip(n4981), .ck(clk), .q(
        \cache_data[14][58] ) );
  dp_1 \cache_data_reg[14][90]  ( .ip(n4949), .ck(clk), .q(
        \cache_data[14][90] ) );
  dp_1 \cache_data_reg[14][122]  ( .ip(n4917), .ck(clk), .q(
        \cache_data[14][122] ) );
  dp_1 \cache_data_reg[15][26]  ( .ip(n4885), .ck(clk), .q(
        \cache_data[15][26] ) );
  dp_1 \cache_data_reg[15][58]  ( .ip(n4853), .ck(clk), .q(
        \cache_data[15][58] ) );
  dp_1 \cache_data_reg[15][90]  ( .ip(n4821), .ck(clk), .q(
        \cache_data[15][90] ) );
  dp_1 \cache_data_reg[15][122]  ( .ip(n4789), .ck(clk), .q(
        \cache_data[15][122] ) );
  dp_1 \iCache_data_wr_reg[27]  ( .ip(n6836), .ck(clk), .q(iCache_data_wr[27])
         );
  dp_1 \cache_data_reg[0][27]  ( .ip(n6804), .ck(clk), .q(\cache_data[0][27] )
         );
  dp_1 \cache_data_reg[0][59]  ( .ip(n6772), .ck(clk), .q(\cache_data[0][59] )
         );
  dp_1 \cache_data_reg[0][91]  ( .ip(n6740), .ck(clk), .q(\cache_data[0][91] )
         );
  dp_1 \cache_data_reg[0][123]  ( .ip(n6708), .ck(clk), .q(
        \cache_data[0][123] ) );
  dp_1 \cache_data_reg[1][27]  ( .ip(n6676), .ck(clk), .q(\cache_data[1][27] )
         );
  dp_1 \cache_data_reg[1][59]  ( .ip(n6644), .ck(clk), .q(\cache_data[1][59] )
         );
  dp_1 \cache_data_reg[1][91]  ( .ip(n6612), .ck(clk), .q(\cache_data[1][91] )
         );
  dp_1 \cache_data_reg[1][123]  ( .ip(n6580), .ck(clk), .q(
        \cache_data[1][123] ) );
  dp_1 \cache_data_reg[2][27]  ( .ip(n6548), .ck(clk), .q(\cache_data[2][27] )
         );
  dp_1 \cache_data_reg[2][59]  ( .ip(n6516), .ck(clk), .q(\cache_data[2][59] )
         );
  dp_1 \cache_data_reg[2][91]  ( .ip(n6484), .ck(clk), .q(\cache_data[2][91] )
         );
  dp_1 \cache_data_reg[2][123]  ( .ip(n6452), .ck(clk), .q(
        \cache_data[2][123] ) );
  dp_1 \cache_data_reg[3][27]  ( .ip(n6420), .ck(clk), .q(\cache_data[3][27] )
         );
  dp_1 \cache_data_reg[3][59]  ( .ip(n6388), .ck(clk), .q(\cache_data[3][59] )
         );
  dp_1 \cache_data_reg[3][91]  ( .ip(n6356), .ck(clk), .q(\cache_data[3][91] )
         );
  dp_1 \cache_data_reg[3][123]  ( .ip(n6324), .ck(clk), .q(
        \cache_data[3][123] ) );
  dp_1 \cache_data_reg[4][27]  ( .ip(n6292), .ck(clk), .q(\cache_data[4][27] )
         );
  dp_1 \cache_data_reg[4][59]  ( .ip(n6260), .ck(clk), .q(\cache_data[4][59] )
         );
  dp_1 \cache_data_reg[4][91]  ( .ip(n6228), .ck(clk), .q(\cache_data[4][91] )
         );
  dp_1 \cache_data_reg[4][123]  ( .ip(n6196), .ck(clk), .q(
        \cache_data[4][123] ) );
  dp_1 \cache_data_reg[5][27]  ( .ip(n6164), .ck(clk), .q(\cache_data[5][27] )
         );
  dp_1 \cache_data_reg[5][59]  ( .ip(n6132), .ck(clk), .q(\cache_data[5][59] )
         );
  dp_1 \cache_data_reg[5][91]  ( .ip(n6100), .ck(clk), .q(\cache_data[5][91] )
         );
  dp_1 \cache_data_reg[5][123]  ( .ip(n6068), .ck(clk), .q(
        \cache_data[5][123] ) );
  dp_1 \cache_data_reg[6][27]  ( .ip(n6036), .ck(clk), .q(\cache_data[6][27] )
         );
  dp_1 \cache_data_reg[6][59]  ( .ip(n6004), .ck(clk), .q(\cache_data[6][59] )
         );
  dp_1 \cache_data_reg[6][91]  ( .ip(n5972), .ck(clk), .q(\cache_data[6][91] )
         );
  dp_1 \cache_data_reg[6][123]  ( .ip(n5940), .ck(clk), .q(
        \cache_data[6][123] ) );
  dp_1 \cache_data_reg[7][27]  ( .ip(n5908), .ck(clk), .q(\cache_data[7][27] )
         );
  dp_1 \cache_data_reg[7][59]  ( .ip(n5876), .ck(clk), .q(\cache_data[7][59] )
         );
  dp_1 \cache_data_reg[7][91]  ( .ip(n5844), .ck(clk), .q(\cache_data[7][91] )
         );
  dp_1 \cache_data_reg[7][123]  ( .ip(n5812), .ck(clk), .q(
        \cache_data[7][123] ) );
  dp_1 \cache_data_reg[8][27]  ( .ip(n5780), .ck(clk), .q(\cache_data[8][27] )
         );
  dp_1 \cache_data_reg[8][59]  ( .ip(n5748), .ck(clk), .q(\cache_data[8][59] )
         );
  dp_1 \cache_data_reg[8][91]  ( .ip(n5716), .ck(clk), .q(\cache_data[8][91] )
         );
  dp_1 \cache_data_reg[8][123]  ( .ip(n5684), .ck(clk), .q(
        \cache_data[8][123] ) );
  dp_1 \cache_data_reg[9][27]  ( .ip(n5652), .ck(clk), .q(\cache_data[9][27] )
         );
  dp_1 \cache_data_reg[9][59]  ( .ip(n5620), .ck(clk), .q(\cache_data[9][59] )
         );
  dp_1 \cache_data_reg[9][91]  ( .ip(n5588), .ck(clk), .q(\cache_data[9][91] )
         );
  dp_1 \cache_data_reg[9][123]  ( .ip(n5556), .ck(clk), .q(
        \cache_data[9][123] ) );
  dp_1 \cache_data_reg[10][27]  ( .ip(n5524), .ck(clk), .q(
        \cache_data[10][27] ) );
  dp_1 \cache_data_reg[10][59]  ( .ip(n5492), .ck(clk), .q(
        \cache_data[10][59] ) );
  dp_1 \cache_data_reg[10][91]  ( .ip(n5460), .ck(clk), .q(
        \cache_data[10][91] ) );
  dp_1 \cache_data_reg[10][123]  ( .ip(n5428), .ck(clk), .q(
        \cache_data[10][123] ) );
  dp_1 \cache_data_reg[11][27]  ( .ip(n5396), .ck(clk), .q(
        \cache_data[11][27] ) );
  dp_1 \cache_data_reg[11][59]  ( .ip(n5364), .ck(clk), .q(
        \cache_data[11][59] ) );
  dp_1 \cache_data_reg[11][91]  ( .ip(n5332), .ck(clk), .q(
        \cache_data[11][91] ) );
  dp_1 \cache_data_reg[11][123]  ( .ip(n5300), .ck(clk), .q(
        \cache_data[11][123] ) );
  dp_1 \cache_data_reg[12][27]  ( .ip(n5268), .ck(clk), .q(
        \cache_data[12][27] ) );
  dp_1 \cache_data_reg[12][59]  ( .ip(n5236), .ck(clk), .q(
        \cache_data[12][59] ) );
  dp_1 \cache_data_reg[12][91]  ( .ip(n5204), .ck(clk), .q(
        \cache_data[12][91] ) );
  dp_1 \cache_data_reg[12][123]  ( .ip(n5172), .ck(clk), .q(
        \cache_data[12][123] ) );
  dp_1 \cache_data_reg[13][27]  ( .ip(n5140), .ck(clk), .q(
        \cache_data[13][27] ) );
  dp_1 \cache_data_reg[13][59]  ( .ip(n5108), .ck(clk), .q(
        \cache_data[13][59] ) );
  dp_1 \cache_data_reg[13][91]  ( .ip(n5076), .ck(clk), .q(
        \cache_data[13][91] ) );
  dp_1 \cache_data_reg[13][123]  ( .ip(n5044), .ck(clk), .q(
        \cache_data[13][123] ) );
  dp_1 \cache_data_reg[14][27]  ( .ip(n5012), .ck(clk), .q(
        \cache_data[14][27] ) );
  dp_1 \cache_data_reg[14][59]  ( .ip(n4980), .ck(clk), .q(
        \cache_data[14][59] ) );
  dp_1 \cache_data_reg[14][91]  ( .ip(n4948), .ck(clk), .q(
        \cache_data[14][91] ) );
  dp_1 \cache_data_reg[14][123]  ( .ip(n4916), .ck(clk), .q(
        \cache_data[14][123] ) );
  dp_1 \cache_data_reg[15][27]  ( .ip(n4884), .ck(clk), .q(
        \cache_data[15][27] ) );
  dp_1 \cache_data_reg[15][59]  ( .ip(n4852), .ck(clk), .q(
        \cache_data[15][59] ) );
  dp_1 \cache_data_reg[15][91]  ( .ip(n4820), .ck(clk), .q(
        \cache_data[15][91] ) );
  dp_1 \cache_data_reg[15][123]  ( .ip(n4788), .ck(clk), .q(
        \cache_data[15][123] ) );
  dp_1 \iCache_data_wr_reg[28]  ( .ip(n6835), .ck(clk), .q(iCache_data_wr[28])
         );
  dp_1 \cache_data_reg[0][28]  ( .ip(n6803), .ck(clk), .q(\cache_data[0][28] )
         );
  dp_1 \cache_data_reg[0][60]  ( .ip(n6771), .ck(clk), .q(\cache_data[0][60] )
         );
  dp_1 \cache_data_reg[0][92]  ( .ip(n6739), .ck(clk), .q(\cache_data[0][92] )
         );
  dp_1 \cache_data_reg[0][124]  ( .ip(n6707), .ck(clk), .q(
        \cache_data[0][124] ) );
  dp_1 \cache_data_reg[1][28]  ( .ip(n6675), .ck(clk), .q(\cache_data[1][28] )
         );
  dp_1 \cache_data_reg[1][60]  ( .ip(n6643), .ck(clk), .q(\cache_data[1][60] )
         );
  dp_1 \cache_data_reg[1][92]  ( .ip(n6611), .ck(clk), .q(\cache_data[1][92] )
         );
  dp_1 \cache_data_reg[1][124]  ( .ip(n6579), .ck(clk), .q(
        \cache_data[1][124] ) );
  dp_1 \cache_data_reg[2][28]  ( .ip(n6547), .ck(clk), .q(\cache_data[2][28] )
         );
  dp_1 \cache_data_reg[2][60]  ( .ip(n6515), .ck(clk), .q(\cache_data[2][60] )
         );
  dp_1 \cache_data_reg[2][92]  ( .ip(n6483), .ck(clk), .q(\cache_data[2][92] )
         );
  dp_1 \cache_data_reg[2][124]  ( .ip(n6451), .ck(clk), .q(
        \cache_data[2][124] ) );
  dp_1 \cache_data_reg[3][28]  ( .ip(n6419), .ck(clk), .q(\cache_data[3][28] )
         );
  dp_1 \cache_data_reg[3][60]  ( .ip(n6387), .ck(clk), .q(\cache_data[3][60] )
         );
  dp_1 \cache_data_reg[3][92]  ( .ip(n6355), .ck(clk), .q(\cache_data[3][92] )
         );
  dp_1 \cache_data_reg[3][124]  ( .ip(n6323), .ck(clk), .q(
        \cache_data[3][124] ) );
  dp_1 \cache_data_reg[4][28]  ( .ip(n6291), .ck(clk), .q(\cache_data[4][28] )
         );
  dp_1 \cache_data_reg[4][60]  ( .ip(n6259), .ck(clk), .q(\cache_data[4][60] )
         );
  dp_1 \cache_data_reg[4][92]  ( .ip(n6227), .ck(clk), .q(\cache_data[4][92] )
         );
  dp_1 \cache_data_reg[4][124]  ( .ip(n6195), .ck(clk), .q(
        \cache_data[4][124] ) );
  dp_1 \cache_data_reg[5][28]  ( .ip(n6163), .ck(clk), .q(\cache_data[5][28] )
         );
  dp_1 \cache_data_reg[5][60]  ( .ip(n6131), .ck(clk), .q(\cache_data[5][60] )
         );
  dp_1 \cache_data_reg[5][92]  ( .ip(n6099), .ck(clk), .q(\cache_data[5][92] )
         );
  dp_1 \cache_data_reg[5][124]  ( .ip(n6067), .ck(clk), .q(
        \cache_data[5][124] ) );
  dp_1 \cache_data_reg[6][28]  ( .ip(n6035), .ck(clk), .q(\cache_data[6][28] )
         );
  dp_1 \cache_data_reg[6][60]  ( .ip(n6003), .ck(clk), .q(\cache_data[6][60] )
         );
  dp_1 \cache_data_reg[6][92]  ( .ip(n5971), .ck(clk), .q(\cache_data[6][92] )
         );
  dp_1 \cache_data_reg[6][124]  ( .ip(n5939), .ck(clk), .q(
        \cache_data[6][124] ) );
  dp_1 \cache_data_reg[7][28]  ( .ip(n5907), .ck(clk), .q(\cache_data[7][28] )
         );
  dp_1 \cache_data_reg[7][60]  ( .ip(n5875), .ck(clk), .q(\cache_data[7][60] )
         );
  dp_1 \cache_data_reg[7][92]  ( .ip(n5843), .ck(clk), .q(\cache_data[7][92] )
         );
  dp_1 \cache_data_reg[7][124]  ( .ip(n5811), .ck(clk), .q(
        \cache_data[7][124] ) );
  dp_1 \cache_data_reg[8][28]  ( .ip(n5779), .ck(clk), .q(\cache_data[8][28] )
         );
  dp_1 \cache_data_reg[8][60]  ( .ip(n5747), .ck(clk), .q(\cache_data[8][60] )
         );
  dp_1 \cache_data_reg[8][92]  ( .ip(n5715), .ck(clk), .q(\cache_data[8][92] )
         );
  dp_1 \cache_data_reg[8][124]  ( .ip(n5683), .ck(clk), .q(
        \cache_data[8][124] ) );
  dp_1 \cache_data_reg[9][28]  ( .ip(n5651), .ck(clk), .q(\cache_data[9][28] )
         );
  dp_1 \cache_data_reg[9][60]  ( .ip(n5619), .ck(clk), .q(\cache_data[9][60] )
         );
  dp_1 \cache_data_reg[9][92]  ( .ip(n5587), .ck(clk), .q(\cache_data[9][92] )
         );
  dp_1 \cache_data_reg[9][124]  ( .ip(n5555), .ck(clk), .q(
        \cache_data[9][124] ) );
  dp_1 \cache_data_reg[10][28]  ( .ip(n5523), .ck(clk), .q(
        \cache_data[10][28] ) );
  dp_1 \cache_data_reg[10][60]  ( .ip(n5491), .ck(clk), .q(
        \cache_data[10][60] ) );
  dp_1 \cache_data_reg[10][92]  ( .ip(n5459), .ck(clk), .q(
        \cache_data[10][92] ) );
  dp_1 \cache_data_reg[10][124]  ( .ip(n5427), .ck(clk), .q(
        \cache_data[10][124] ) );
  dp_1 \cache_data_reg[11][28]  ( .ip(n5395), .ck(clk), .q(
        \cache_data[11][28] ) );
  dp_1 \cache_data_reg[11][60]  ( .ip(n5363), .ck(clk), .q(
        \cache_data[11][60] ) );
  dp_1 \cache_data_reg[11][92]  ( .ip(n5331), .ck(clk), .q(
        \cache_data[11][92] ) );
  dp_1 \cache_data_reg[11][124]  ( .ip(n5299), .ck(clk), .q(
        \cache_data[11][124] ) );
  dp_1 \cache_data_reg[12][28]  ( .ip(n5267), .ck(clk), .q(
        \cache_data[12][28] ) );
  dp_1 \cache_data_reg[12][60]  ( .ip(n5235), .ck(clk), .q(
        \cache_data[12][60] ) );
  dp_1 \cache_data_reg[12][92]  ( .ip(n5203), .ck(clk), .q(
        \cache_data[12][92] ) );
  dp_1 \cache_data_reg[12][124]  ( .ip(n5171), .ck(clk), .q(
        \cache_data[12][124] ) );
  dp_1 \cache_data_reg[13][28]  ( .ip(n5139), .ck(clk), .q(
        \cache_data[13][28] ) );
  dp_1 \cache_data_reg[13][60]  ( .ip(n5107), .ck(clk), .q(
        \cache_data[13][60] ) );
  dp_1 \cache_data_reg[13][92]  ( .ip(n5075), .ck(clk), .q(
        \cache_data[13][92] ) );
  dp_1 \cache_data_reg[13][124]  ( .ip(n5043), .ck(clk), .q(
        \cache_data[13][124] ) );
  dp_1 \cache_data_reg[14][28]  ( .ip(n5011), .ck(clk), .q(
        \cache_data[14][28] ) );
  dp_1 \cache_data_reg[14][60]  ( .ip(n4979), .ck(clk), .q(
        \cache_data[14][60] ) );
  dp_1 \cache_data_reg[14][92]  ( .ip(n4947), .ck(clk), .q(
        \cache_data[14][92] ) );
  dp_1 \cache_data_reg[14][124]  ( .ip(n4915), .ck(clk), .q(
        \cache_data[14][124] ) );
  dp_1 \cache_data_reg[15][28]  ( .ip(n4883), .ck(clk), .q(
        \cache_data[15][28] ) );
  dp_1 \cache_data_reg[15][60]  ( .ip(n4851), .ck(clk), .q(
        \cache_data[15][60] ) );
  dp_1 \cache_data_reg[15][92]  ( .ip(n4819), .ck(clk), .q(
        \cache_data[15][92] ) );
  dp_1 \cache_data_reg[15][124]  ( .ip(n4787), .ck(clk), .q(
        \cache_data[15][124] ) );
  dp_1 \iCache_data_wr_reg[29]  ( .ip(n6834), .ck(clk), .q(iCache_data_wr[29])
         );
  dp_1 \cache_data_reg[0][29]  ( .ip(n6802), .ck(clk), .q(\cache_data[0][29] )
         );
  dp_1 \cache_data_reg[0][61]  ( .ip(n6770), .ck(clk), .q(\cache_data[0][61] )
         );
  dp_1 \cache_data_reg[0][93]  ( .ip(n6738), .ck(clk), .q(\cache_data[0][93] )
         );
  dp_1 \cache_data_reg[0][125]  ( .ip(n6706), .ck(clk), .q(
        \cache_data[0][125] ) );
  dp_1 \cache_data_reg[1][29]  ( .ip(n6674), .ck(clk), .q(\cache_data[1][29] )
         );
  dp_1 \cache_data_reg[1][61]  ( .ip(n6642), .ck(clk), .q(\cache_data[1][61] )
         );
  dp_1 \cache_data_reg[1][93]  ( .ip(n6610), .ck(clk), .q(\cache_data[1][93] )
         );
  dp_1 \cache_data_reg[1][125]  ( .ip(n6578), .ck(clk), .q(
        \cache_data[1][125] ) );
  dp_1 \cache_data_reg[2][29]  ( .ip(n6546), .ck(clk), .q(\cache_data[2][29] )
         );
  dp_1 \cache_data_reg[2][61]  ( .ip(n6514), .ck(clk), .q(\cache_data[2][61] )
         );
  dp_1 \cache_data_reg[2][93]  ( .ip(n6482), .ck(clk), .q(\cache_data[2][93] )
         );
  dp_1 \cache_data_reg[2][125]  ( .ip(n6450), .ck(clk), .q(
        \cache_data[2][125] ) );
  dp_1 \cache_data_reg[3][29]  ( .ip(n6418), .ck(clk), .q(\cache_data[3][29] )
         );
  dp_1 \cache_data_reg[3][61]  ( .ip(n6386), .ck(clk), .q(\cache_data[3][61] )
         );
  dp_1 \cache_data_reg[3][93]  ( .ip(n6354), .ck(clk), .q(\cache_data[3][93] )
         );
  dp_1 \cache_data_reg[3][125]  ( .ip(n6322), .ck(clk), .q(
        \cache_data[3][125] ) );
  dp_1 \cache_data_reg[4][29]  ( .ip(n6290), .ck(clk), .q(\cache_data[4][29] )
         );
  dp_1 \cache_data_reg[4][61]  ( .ip(n6258), .ck(clk), .q(\cache_data[4][61] )
         );
  dp_1 \cache_data_reg[4][93]  ( .ip(n6226), .ck(clk), .q(\cache_data[4][93] )
         );
  dp_1 \cache_data_reg[4][125]  ( .ip(n6194), .ck(clk), .q(
        \cache_data[4][125] ) );
  dp_1 \cache_data_reg[5][29]  ( .ip(n6162), .ck(clk), .q(\cache_data[5][29] )
         );
  dp_1 \cache_data_reg[5][61]  ( .ip(n6130), .ck(clk), .q(\cache_data[5][61] )
         );
  dp_1 \cache_data_reg[5][93]  ( .ip(n6098), .ck(clk), .q(\cache_data[5][93] )
         );
  dp_1 \cache_data_reg[5][125]  ( .ip(n6066), .ck(clk), .q(
        \cache_data[5][125] ) );
  dp_1 \cache_data_reg[6][29]  ( .ip(n6034), .ck(clk), .q(\cache_data[6][29] )
         );
  dp_1 \cache_data_reg[6][61]  ( .ip(n6002), .ck(clk), .q(\cache_data[6][61] )
         );
  dp_1 \cache_data_reg[6][93]  ( .ip(n5970), .ck(clk), .q(\cache_data[6][93] )
         );
  dp_1 \cache_data_reg[6][125]  ( .ip(n5938), .ck(clk), .q(
        \cache_data[6][125] ) );
  dp_1 \cache_data_reg[7][29]  ( .ip(n5906), .ck(clk), .q(\cache_data[7][29] )
         );
  dp_1 \cache_data_reg[7][61]  ( .ip(n5874), .ck(clk), .q(\cache_data[7][61] )
         );
  dp_1 \cache_data_reg[7][93]  ( .ip(n5842), .ck(clk), .q(\cache_data[7][93] )
         );
  dp_1 \cache_data_reg[7][125]  ( .ip(n5810), .ck(clk), .q(
        \cache_data[7][125] ) );
  dp_1 \cache_data_reg[8][29]  ( .ip(n5778), .ck(clk), .q(\cache_data[8][29] )
         );
  dp_1 \cache_data_reg[8][61]  ( .ip(n5746), .ck(clk), .q(\cache_data[8][61] )
         );
  dp_1 \cache_data_reg[8][93]  ( .ip(n5714), .ck(clk), .q(\cache_data[8][93] )
         );
  dp_1 \cache_data_reg[8][125]  ( .ip(n5682), .ck(clk), .q(
        \cache_data[8][125] ) );
  dp_1 \cache_data_reg[9][29]  ( .ip(n5650), .ck(clk), .q(\cache_data[9][29] )
         );
  dp_1 \cache_data_reg[9][61]  ( .ip(n5618), .ck(clk), .q(\cache_data[9][61] )
         );
  dp_1 \cache_data_reg[9][93]  ( .ip(n5586), .ck(clk), .q(\cache_data[9][93] )
         );
  dp_1 \cache_data_reg[9][125]  ( .ip(n5554), .ck(clk), .q(
        \cache_data[9][125] ) );
  dp_1 \cache_data_reg[10][29]  ( .ip(n5522), .ck(clk), .q(
        \cache_data[10][29] ) );
  dp_1 \cache_data_reg[10][61]  ( .ip(n5490), .ck(clk), .q(
        \cache_data[10][61] ) );
  dp_1 \cache_data_reg[10][93]  ( .ip(n5458), .ck(clk), .q(
        \cache_data[10][93] ) );
  dp_1 \cache_data_reg[10][125]  ( .ip(n5426), .ck(clk), .q(
        \cache_data[10][125] ) );
  dp_1 \cache_data_reg[11][29]  ( .ip(n5394), .ck(clk), .q(
        \cache_data[11][29] ) );
  dp_1 \cache_data_reg[11][61]  ( .ip(n5362), .ck(clk), .q(
        \cache_data[11][61] ) );
  dp_1 \cache_data_reg[11][93]  ( .ip(n5330), .ck(clk), .q(
        \cache_data[11][93] ) );
  dp_1 \cache_data_reg[11][125]  ( .ip(n5298), .ck(clk), .q(
        \cache_data[11][125] ) );
  dp_1 \cache_data_reg[12][29]  ( .ip(n5266), .ck(clk), .q(
        \cache_data[12][29] ) );
  dp_1 \cache_data_reg[12][61]  ( .ip(n5234), .ck(clk), .q(
        \cache_data[12][61] ) );
  dp_1 \cache_data_reg[12][93]  ( .ip(n5202), .ck(clk), .q(
        \cache_data[12][93] ) );
  dp_1 \cache_data_reg[12][125]  ( .ip(n5170), .ck(clk), .q(
        \cache_data[12][125] ) );
  dp_1 \cache_data_reg[13][29]  ( .ip(n5138), .ck(clk), .q(
        \cache_data[13][29] ) );
  dp_1 \cache_data_reg[13][61]  ( .ip(n5106), .ck(clk), .q(
        \cache_data[13][61] ) );
  dp_1 \cache_data_reg[13][93]  ( .ip(n5074), .ck(clk), .q(
        \cache_data[13][93] ) );
  dp_1 \cache_data_reg[13][125]  ( .ip(n5042), .ck(clk), .q(
        \cache_data[13][125] ) );
  dp_1 \cache_data_reg[14][29]  ( .ip(n5010), .ck(clk), .q(
        \cache_data[14][29] ) );
  dp_1 \cache_data_reg[14][61]  ( .ip(n4978), .ck(clk), .q(
        \cache_data[14][61] ) );
  dp_1 \cache_data_reg[14][93]  ( .ip(n4946), .ck(clk), .q(
        \cache_data[14][93] ) );
  dp_1 \cache_data_reg[14][125]  ( .ip(n4914), .ck(clk), .q(
        \cache_data[14][125] ) );
  dp_1 \cache_data_reg[15][29]  ( .ip(n4882), .ck(clk), .q(
        \cache_data[15][29] ) );
  dp_1 \cache_data_reg[15][61]  ( .ip(n4850), .ck(clk), .q(
        \cache_data[15][61] ) );
  dp_1 \cache_data_reg[15][93]  ( .ip(n4818), .ck(clk), .q(
        \cache_data[15][93] ) );
  dp_1 \cache_data_reg[15][125]  ( .ip(n4786), .ck(clk), .q(
        \cache_data[15][125] ) );
  dp_1 \iCache_data_wr_reg[30]  ( .ip(n6833), .ck(clk), .q(iCache_data_wr[30])
         );
  dp_1 \cache_data_reg[0][30]  ( .ip(n6801), .ck(clk), .q(\cache_data[0][30] )
         );
  dp_1 \cache_data_reg[0][62]  ( .ip(n6769), .ck(clk), .q(\cache_data[0][62] )
         );
  dp_1 \cache_data_reg[0][94]  ( .ip(n6737), .ck(clk), .q(\cache_data[0][94] )
         );
  dp_1 \cache_data_reg[0][126]  ( .ip(n6705), .ck(clk), .q(
        \cache_data[0][126] ) );
  dp_1 \cache_data_reg[1][30]  ( .ip(n6673), .ck(clk), .q(\cache_data[1][30] )
         );
  dp_1 \cache_data_reg[1][62]  ( .ip(n6641), .ck(clk), .q(\cache_data[1][62] )
         );
  dp_1 \cache_data_reg[1][94]  ( .ip(n6609), .ck(clk), .q(\cache_data[1][94] )
         );
  dp_1 \cache_data_reg[1][126]  ( .ip(n6577), .ck(clk), .q(
        \cache_data[1][126] ) );
  dp_1 \cache_data_reg[2][30]  ( .ip(n6545), .ck(clk), .q(\cache_data[2][30] )
         );
  dp_1 \cache_data_reg[2][62]  ( .ip(n6513), .ck(clk), .q(\cache_data[2][62] )
         );
  dp_1 \cache_data_reg[2][94]  ( .ip(n6481), .ck(clk), .q(\cache_data[2][94] )
         );
  dp_1 \cache_data_reg[2][126]  ( .ip(n6449), .ck(clk), .q(
        \cache_data[2][126] ) );
  dp_1 \cache_data_reg[3][30]  ( .ip(n6417), .ck(clk), .q(\cache_data[3][30] )
         );
  dp_1 \cache_data_reg[3][62]  ( .ip(n6385), .ck(clk), .q(\cache_data[3][62] )
         );
  dp_1 \cache_data_reg[3][94]  ( .ip(n6353), .ck(clk), .q(\cache_data[3][94] )
         );
  dp_1 \cache_data_reg[3][126]  ( .ip(n6321), .ck(clk), .q(
        \cache_data[3][126] ) );
  dp_1 \cache_data_reg[4][30]  ( .ip(n6289), .ck(clk), .q(\cache_data[4][30] )
         );
  dp_1 \cache_data_reg[4][62]  ( .ip(n6257), .ck(clk), .q(\cache_data[4][62] )
         );
  dp_1 \cache_data_reg[4][94]  ( .ip(n6225), .ck(clk), .q(\cache_data[4][94] )
         );
  dp_1 \cache_data_reg[4][126]  ( .ip(n6193), .ck(clk), .q(
        \cache_data[4][126] ) );
  dp_1 \cache_data_reg[5][30]  ( .ip(n6161), .ck(clk), .q(\cache_data[5][30] )
         );
  dp_1 \cache_data_reg[5][62]  ( .ip(n6129), .ck(clk), .q(\cache_data[5][62] )
         );
  dp_1 \cache_data_reg[5][94]  ( .ip(n6097), .ck(clk), .q(\cache_data[5][94] )
         );
  dp_1 \cache_data_reg[5][126]  ( .ip(n6065), .ck(clk), .q(
        \cache_data[5][126] ) );
  dp_1 \cache_data_reg[6][30]  ( .ip(n6033), .ck(clk), .q(\cache_data[6][30] )
         );
  dp_1 \cache_data_reg[6][62]  ( .ip(n6001), .ck(clk), .q(\cache_data[6][62] )
         );
  dp_1 \cache_data_reg[6][94]  ( .ip(n5969), .ck(clk), .q(\cache_data[6][94] )
         );
  dp_1 \cache_data_reg[6][126]  ( .ip(n5937), .ck(clk), .q(
        \cache_data[6][126] ) );
  dp_1 \cache_data_reg[7][30]  ( .ip(n5905), .ck(clk), .q(\cache_data[7][30] )
         );
  dp_1 \cache_data_reg[7][62]  ( .ip(n5873), .ck(clk), .q(\cache_data[7][62] )
         );
  dp_1 \cache_data_reg[7][94]  ( .ip(n5841), .ck(clk), .q(\cache_data[7][94] )
         );
  dp_1 \cache_data_reg[7][126]  ( .ip(n5809), .ck(clk), .q(
        \cache_data[7][126] ) );
  dp_1 \cache_data_reg[8][30]  ( .ip(n5777), .ck(clk), .q(\cache_data[8][30] )
         );
  dp_1 \cache_data_reg[8][62]  ( .ip(n5745), .ck(clk), .q(\cache_data[8][62] )
         );
  dp_1 \cache_data_reg[8][94]  ( .ip(n5713), .ck(clk), .q(\cache_data[8][94] )
         );
  dp_1 \cache_data_reg[8][126]  ( .ip(n5681), .ck(clk), .q(
        \cache_data[8][126] ) );
  dp_1 \cache_data_reg[9][30]  ( .ip(n5649), .ck(clk), .q(\cache_data[9][30] )
         );
  dp_1 \cache_data_reg[9][62]  ( .ip(n5617), .ck(clk), .q(\cache_data[9][62] )
         );
  dp_1 \cache_data_reg[9][94]  ( .ip(n5585), .ck(clk), .q(\cache_data[9][94] )
         );
  dp_1 \cache_data_reg[9][126]  ( .ip(n5553), .ck(clk), .q(
        \cache_data[9][126] ) );
  dp_1 \cache_data_reg[10][30]  ( .ip(n5521), .ck(clk), .q(
        \cache_data[10][30] ) );
  dp_1 \cache_data_reg[10][62]  ( .ip(n5489), .ck(clk), .q(
        \cache_data[10][62] ) );
  dp_1 \cache_data_reg[10][94]  ( .ip(n5457), .ck(clk), .q(
        \cache_data[10][94] ) );
  dp_1 \cache_data_reg[10][126]  ( .ip(n5425), .ck(clk), .q(
        \cache_data[10][126] ) );
  dp_1 \cache_data_reg[11][30]  ( .ip(n5393), .ck(clk), .q(
        \cache_data[11][30] ) );
  dp_1 \cache_data_reg[11][62]  ( .ip(n5361), .ck(clk), .q(
        \cache_data[11][62] ) );
  dp_1 \cache_data_reg[11][94]  ( .ip(n5329), .ck(clk), .q(
        \cache_data[11][94] ) );
  dp_1 \cache_data_reg[11][126]  ( .ip(n5297), .ck(clk), .q(
        \cache_data[11][126] ) );
  dp_1 \cache_data_reg[12][30]  ( .ip(n5265), .ck(clk), .q(
        \cache_data[12][30] ) );
  dp_1 \cache_data_reg[12][62]  ( .ip(n5233), .ck(clk), .q(
        \cache_data[12][62] ) );
  dp_1 \cache_data_reg[12][94]  ( .ip(n5201), .ck(clk), .q(
        \cache_data[12][94] ) );
  dp_1 \cache_data_reg[12][126]  ( .ip(n5169), .ck(clk), .q(
        \cache_data[12][126] ) );
  dp_1 \cache_data_reg[13][30]  ( .ip(n5137), .ck(clk), .q(
        \cache_data[13][30] ) );
  dp_1 \cache_data_reg[13][62]  ( .ip(n5105), .ck(clk), .q(
        \cache_data[13][62] ) );
  dp_1 \cache_data_reg[13][94]  ( .ip(n5073), .ck(clk), .q(
        \cache_data[13][94] ) );
  dp_1 \cache_data_reg[13][126]  ( .ip(n5041), .ck(clk), .q(
        \cache_data[13][126] ) );
  dp_1 \cache_data_reg[14][30]  ( .ip(n5009), .ck(clk), .q(
        \cache_data[14][30] ) );
  dp_1 \cache_data_reg[14][62]  ( .ip(n4977), .ck(clk), .q(
        \cache_data[14][62] ) );
  dp_1 \cache_data_reg[14][94]  ( .ip(n4945), .ck(clk), .q(
        \cache_data[14][94] ) );
  dp_1 \cache_data_reg[14][126]  ( .ip(n4913), .ck(clk), .q(
        \cache_data[14][126] ) );
  dp_1 \cache_data_reg[15][30]  ( .ip(n4881), .ck(clk), .q(
        \cache_data[15][30] ) );
  dp_1 \cache_data_reg[15][62]  ( .ip(n4849), .ck(clk), .q(
        \cache_data[15][62] ) );
  dp_1 \cache_data_reg[15][94]  ( .ip(n4817), .ck(clk), .q(
        \cache_data[15][94] ) );
  dp_1 \cache_data_reg[15][126]  ( .ip(n4785), .ck(clk), .q(
        \cache_data[15][126] ) );
  dp_1 \iCache_data_wr_reg[31]  ( .ip(n6832), .ck(clk), .q(iCache_data_wr[31])
         );
  dp_1 \cache_data_reg[0][31]  ( .ip(n6800), .ck(clk), .q(\cache_data[0][31] )
         );
  dp_1 \cache_data_reg[0][63]  ( .ip(n6768), .ck(clk), .q(\cache_data[0][63] )
         );
  dp_1 \cache_data_reg[0][95]  ( .ip(n6736), .ck(clk), .q(\cache_data[0][95] )
         );
  dp_1 \cache_data_reg[0][127]  ( .ip(n6704), .ck(clk), .q(
        \cache_data[0][127] ) );
  dp_1 \cache_data_reg[1][31]  ( .ip(n6672), .ck(clk), .q(\cache_data[1][31] )
         );
  dp_1 \cache_data_reg[1][63]  ( .ip(n6640), .ck(clk), .q(\cache_data[1][63] )
         );
  dp_1 \cache_data_reg[1][95]  ( .ip(n6608), .ck(clk), .q(\cache_data[1][95] )
         );
  dp_1 \cache_data_reg[1][127]  ( .ip(n6576), .ck(clk), .q(
        \cache_data[1][127] ) );
  dp_1 \cache_data_reg[2][31]  ( .ip(n6544), .ck(clk), .q(\cache_data[2][31] )
         );
  dp_1 \cache_data_reg[2][63]  ( .ip(n6512), .ck(clk), .q(\cache_data[2][63] )
         );
  dp_1 \cache_data_reg[2][95]  ( .ip(n6480), .ck(clk), .q(\cache_data[2][95] )
         );
  dp_1 \cache_data_reg[2][127]  ( .ip(n6448), .ck(clk), .q(
        \cache_data[2][127] ) );
  dp_1 \cache_data_reg[3][31]  ( .ip(n6416), .ck(clk), .q(\cache_data[3][31] )
         );
  dp_1 \cache_data_reg[3][63]  ( .ip(n6384), .ck(clk), .q(\cache_data[3][63] )
         );
  dp_1 \cache_data_reg[3][95]  ( .ip(n6352), .ck(clk), .q(\cache_data[3][95] )
         );
  dp_1 \cache_data_reg[3][127]  ( .ip(n6320), .ck(clk), .q(
        \cache_data[3][127] ) );
  dp_1 \cache_data_reg[4][31]  ( .ip(n6288), .ck(clk), .q(\cache_data[4][31] )
         );
  dp_1 \cache_data_reg[4][63]  ( .ip(n6256), .ck(clk), .q(\cache_data[4][63] )
         );
  dp_1 \cache_data_reg[4][95]  ( .ip(n6224), .ck(clk), .q(\cache_data[4][95] )
         );
  dp_1 \cache_data_reg[4][127]  ( .ip(n6192), .ck(clk), .q(
        \cache_data[4][127] ) );
  dp_1 \cache_data_reg[5][31]  ( .ip(n6160), .ck(clk), .q(\cache_data[5][31] )
         );
  dp_1 \cache_data_reg[5][63]  ( .ip(n6128), .ck(clk), .q(\cache_data[5][63] )
         );
  dp_1 \cache_data_reg[5][95]  ( .ip(n6096), .ck(clk), .q(\cache_data[5][95] )
         );
  dp_1 \cache_data_reg[5][127]  ( .ip(n6064), .ck(clk), .q(
        \cache_data[5][127] ) );
  dp_1 \cache_data_reg[6][31]  ( .ip(n6032), .ck(clk), .q(\cache_data[6][31] )
         );
  dp_1 \cache_data_reg[6][63]  ( .ip(n6000), .ck(clk), .q(\cache_data[6][63] )
         );
  dp_1 \cache_data_reg[6][95]  ( .ip(n5968), .ck(clk), .q(\cache_data[6][95] )
         );
  dp_1 \cache_data_reg[6][127]  ( .ip(n5936), .ck(clk), .q(
        \cache_data[6][127] ) );
  dp_1 \cache_data_reg[7][31]  ( .ip(n5904), .ck(clk), .q(\cache_data[7][31] )
         );
  dp_1 \cache_data_reg[7][63]  ( .ip(n5872), .ck(clk), .q(\cache_data[7][63] )
         );
  dp_1 \cache_data_reg[7][95]  ( .ip(n5840), .ck(clk), .q(\cache_data[7][95] )
         );
  dp_1 \cache_data_reg[7][127]  ( .ip(n5808), .ck(clk), .q(
        \cache_data[7][127] ) );
  dp_1 \cache_data_reg[8][31]  ( .ip(n5776), .ck(clk), .q(\cache_data[8][31] )
         );
  dp_1 \cache_data_reg[8][63]  ( .ip(n5744), .ck(clk), .q(\cache_data[8][63] )
         );
  dp_1 \cache_data_reg[8][95]  ( .ip(n5712), .ck(clk), .q(\cache_data[8][95] )
         );
  dp_1 \cache_data_reg[8][127]  ( .ip(n5680), .ck(clk), .q(
        \cache_data[8][127] ) );
  dp_1 \cache_data_reg[9][31]  ( .ip(n5648), .ck(clk), .q(\cache_data[9][31] )
         );
  dp_1 \cache_data_reg[9][63]  ( .ip(n5616), .ck(clk), .q(\cache_data[9][63] )
         );
  dp_1 \cache_data_reg[9][95]  ( .ip(n5584), .ck(clk), .q(\cache_data[9][95] )
         );
  dp_1 \cache_data_reg[9][127]  ( .ip(n5552), .ck(clk), .q(
        \cache_data[9][127] ) );
  dp_1 \cache_data_reg[10][31]  ( .ip(n5520), .ck(clk), .q(
        \cache_data[10][31] ) );
  dp_1 \cache_data_reg[10][63]  ( .ip(n5488), .ck(clk), .q(
        \cache_data[10][63] ) );
  dp_1 \cache_data_reg[10][95]  ( .ip(n5456), .ck(clk), .q(
        \cache_data[10][95] ) );
  dp_1 \cache_data_reg[10][127]  ( .ip(n5424), .ck(clk), .q(
        \cache_data[10][127] ) );
  dp_1 \cache_data_reg[11][31]  ( .ip(n5392), .ck(clk), .q(
        \cache_data[11][31] ) );
  dp_1 \cache_data_reg[11][63]  ( .ip(n5360), .ck(clk), .q(
        \cache_data[11][63] ) );
  dp_1 \cache_data_reg[11][95]  ( .ip(n5328), .ck(clk), .q(
        \cache_data[11][95] ) );
  dp_1 \cache_data_reg[11][127]  ( .ip(n5296), .ck(clk), .q(
        \cache_data[11][127] ) );
  dp_1 \cache_data_reg[12][31]  ( .ip(n5264), .ck(clk), .q(
        \cache_data[12][31] ) );
  dp_1 \cache_data_reg[12][63]  ( .ip(n5232), .ck(clk), .q(
        \cache_data[12][63] ) );
  dp_1 \cache_data_reg[12][95]  ( .ip(n5200), .ck(clk), .q(
        \cache_data[12][95] ) );
  dp_1 \cache_data_reg[12][127]  ( .ip(n5168), .ck(clk), .q(
        \cache_data[12][127] ) );
  dp_1 \cache_data_reg[13][31]  ( .ip(n5136), .ck(clk), .q(
        \cache_data[13][31] ) );
  dp_1 \cache_data_reg[13][63]  ( .ip(n5104), .ck(clk), .q(
        \cache_data[13][63] ) );
  dp_1 \cache_data_reg[13][95]  ( .ip(n5072), .ck(clk), .q(
        \cache_data[13][95] ) );
  dp_1 \cache_data_reg[13][127]  ( .ip(n5040), .ck(clk), .q(
        \cache_data[13][127] ) );
  dp_1 \cache_data_reg[14][31]  ( .ip(n5008), .ck(clk), .q(
        \cache_data[14][31] ) );
  dp_1 \cache_data_reg[14][63]  ( .ip(n4976), .ck(clk), .q(
        \cache_data[14][63] ) );
  dp_1 \cache_data_reg[14][95]  ( .ip(n4944), .ck(clk), .q(
        \cache_data[14][95] ) );
  dp_1 \cache_data_reg[14][127]  ( .ip(n4912), .ck(clk), .q(
        \cache_data[14][127] ) );
  dp_1 \cache_data_reg[15][31]  ( .ip(n4880), .ck(clk), .q(
        \cache_data[15][31] ) );
  dp_1 \cache_data_reg[15][63]  ( .ip(n4848), .ck(clk), .q(
        \cache_data[15][63] ) );
  dp_1 \cache_data_reg[15][95]  ( .ip(n4816), .ck(clk), .q(
        \cache_data[15][95] ) );
  dp_1 \cache_data_reg[15][127]  ( .ip(n4784), .ck(clk), .q(
        \cache_data[15][127] ) );
  drp_1 \cache_miss_count_reg[31]  ( .ip(n4750), .ck(clk), .rb(n12330), .q(
        cache_miss_count[31]) );
  drp_1 \cache_miss_count_reg[30]  ( .ip(n4749), .ck(clk), .rb(n12330), .q(
        cache_miss_count[30]) );
  drp_1 \cache_miss_count_reg[29]  ( .ip(n4748), .ck(clk), .rb(n12330), .q(
        cache_miss_count[29]) );
  drp_1 \cache_miss_count_reg[28]  ( .ip(n4747), .ck(clk), .rb(n12330), .q(
        cache_miss_count[28]) );
  drp_1 \cache_miss_count_reg[27]  ( .ip(n4746), .ck(clk), .rb(n12329), .q(
        cache_miss_count[27]) );
  drp_1 \cache_miss_count_reg[26]  ( .ip(n4745), .ck(clk), .rb(n12329), .q(
        cache_miss_count[26]) );
  drp_1 \cache_miss_count_reg[25]  ( .ip(n4744), .ck(clk), .rb(n12329), .q(
        cache_miss_count[25]) );
  drp_1 \cache_miss_count_reg[24]  ( .ip(n4743), .ck(clk), .rb(n12329), .q(
        cache_miss_count[24]) );
  drp_1 \cache_miss_count_reg[23]  ( .ip(n4742), .ck(clk), .rb(n12329), .q(
        cache_miss_count[23]) );
  drp_1 \cache_miss_count_reg[22]  ( .ip(n4741), .ck(clk), .rb(n12329), .q(
        cache_miss_count[22]) );
  drp_1 \cache_miss_count_reg[21]  ( .ip(n4740), .ck(clk), .rb(n12329), .q(
        cache_miss_count[21]) );
  drp_1 \cache_miss_count_reg[20]  ( .ip(n4739), .ck(clk), .rb(n12329), .q(
        cache_miss_count[20]) );
  drp_1 \cache_miss_count_reg[19]  ( .ip(n4738), .ck(clk), .rb(n12329), .q(
        cache_miss_count[19]) );
  drp_1 \cache_miss_count_reg[18]  ( .ip(n4737), .ck(clk), .rb(n12329), .q(
        cache_miss_count[18]) );
  drp_1 \cache_miss_count_reg[17]  ( .ip(n4736), .ck(clk), .rb(n12329), .q(
        cache_miss_count[17]) );
  drp_1 \cache_miss_count_reg[16]  ( .ip(n4735), .ck(clk), .rb(n12329), .q(
        cache_miss_count[16]) );
  drp_1 \cache_miss_count_reg[15]  ( .ip(n4734), .ck(clk), .rb(n12326), .q(
        cache_miss_count[15]) );
  drp_1 \cache_miss_count_reg[14]  ( .ip(n4733), .ck(clk), .rb(n12322), .q(
        cache_miss_count[14]) );
  drp_1 \cache_miss_count_reg[13]  ( .ip(n4732), .ck(clk), .rb(n12322), .q(
        cache_miss_count[13]) );
  drp_1 \cache_miss_count_reg[12]  ( .ip(n4731), .ck(clk), .rb(n12322), .q(
        cache_miss_count[12]) );
  drp_1 \cache_miss_count_reg[11]  ( .ip(n4730), .ck(clk), .rb(n12322), .q(
        cache_miss_count[11]) );
  drp_1 \cache_miss_count_reg[10]  ( .ip(n4729), .ck(clk), .rb(n12322), .q(
        cache_miss_count[10]) );
  drp_1 \cache_miss_count_reg[9]  ( .ip(n4728), .ck(clk), .rb(n12322), .q(
        cache_miss_count[9]) );
  drp_1 \cache_miss_count_reg[8]  ( .ip(n4727), .ck(clk), .rb(n12322), .q(
        cache_miss_count[8]) );
  drp_1 \cache_miss_count_reg[7]  ( .ip(n4726), .ck(clk), .rb(n12322), .q(
        cache_miss_count[7]) );
  drp_1 \cache_miss_count_reg[6]  ( .ip(n4725), .ck(clk), .rb(n12322), .q(
        cache_miss_count[6]) );
  drp_1 \cache_miss_count_reg[5]  ( .ip(n4724), .ck(clk), .rb(n12322), .q(
        cache_miss_count[5]) );
  drp_1 \cache_miss_count_reg[4]  ( .ip(n4723), .ck(clk), .rb(n12322), .q(
        cache_miss_count[4]) );
  drp_1 \cache_miss_count_reg[3]  ( .ip(n4722), .ck(clk), .rb(n12328), .q(
        cache_miss_count[3]) );
  drp_1 \cache_miss_count_reg[2]  ( .ip(n4721), .ck(clk), .rb(n12328), .q(
        cache_miss_count[2]) );
  drp_1 \cache_miss_count_reg[1]  ( .ip(n4720), .ck(clk), .rb(n12328), .q(
        cache_miss_count[1]) );
  drp_1 \cache_miss_count_reg[0]  ( .ip(n4719), .ck(clk), .rb(n12328), .q(
        cache_miss_count[0]) );
  drp_1 \cache_hit_count_reg[31]  ( .ip(n4718), .ck(clk), .rb(n12328), .q(
        cache_hit_count[31]) );
  drp_1 \cache_hit_count_reg[30]  ( .ip(n4717), .ck(clk), .rb(n12328), .q(
        cache_hit_count[30]) );
  drp_1 \cache_hit_count_reg[29]  ( .ip(n4716), .ck(clk), .rb(n12328), .q(
        cache_hit_count[29]) );
  drp_1 \cache_hit_count_reg[28]  ( .ip(n4715), .ck(clk), .rb(n12328), .q(
        cache_hit_count[28]) );
  drp_1 \cache_hit_count_reg[27]  ( .ip(n4714), .ck(clk), .rb(n12328), .q(
        cache_hit_count[27]) );
  drp_1 \cache_hit_count_reg[26]  ( .ip(n4713), .ck(clk), .rb(n12328), .q(
        cache_hit_count[26]) );
  drp_1 \cache_hit_count_reg[25]  ( .ip(n4712), .ck(clk), .rb(n12328), .q(
        cache_hit_count[25]) );
  drp_1 \cache_hit_count_reg[24]  ( .ip(n4711), .ck(clk), .rb(n12328), .q(
        cache_hit_count[24]) );
  drp_1 \cache_hit_count_reg[23]  ( .ip(n4710), .ck(clk), .rb(n12333), .q(
        cache_hit_count[23]) );
  drp_1 \cache_hit_count_reg[22]  ( .ip(n4709), .ck(clk), .rb(n12333), .q(
        cache_hit_count[22]) );
  drp_1 \cache_hit_count_reg[21]  ( .ip(n4708), .ck(clk), .rb(n12333), .q(
        cache_hit_count[21]) );
  drp_1 \cache_hit_count_reg[20]  ( .ip(n4707), .ck(clk), .rb(n12333), .q(
        cache_hit_count[20]) );
  drp_1 \cache_hit_count_reg[19]  ( .ip(n4706), .ck(clk), .rb(n12322), .q(
        cache_hit_count[19]) );
  drp_1 \cache_hit_count_reg[18]  ( .ip(n4705), .ck(clk), .rb(n12322), .q(
        cache_hit_count[18]) );
  drp_1 \cache_hit_count_reg[17]  ( .ip(n4704), .ck(clk), .rb(n12322), .q(
        cache_hit_count[17]) );
  drp_1 \cache_hit_count_reg[16]  ( .ip(n4703), .ck(clk), .rb(n12322), .q(
        cache_hit_count[16]) );
  drp_1 \cache_hit_count_reg[15]  ( .ip(n4702), .ck(clk), .rb(n12326), .q(
        cache_hit_count[15]) );
  drp_1 \cache_hit_count_reg[14]  ( .ip(n4701), .ck(clk), .rb(n12326), .q(
        cache_hit_count[14]) );
  drp_1 \cache_hit_count_reg[13]  ( .ip(n4700), .ck(clk), .rb(n12326), .q(
        cache_hit_count[13]) );
  drp_1 \cache_hit_count_reg[12]  ( .ip(n4699), .ck(clk), .rb(n12326), .q(
        cache_hit_count[12]) );
  drp_1 \cache_hit_count_reg[11]  ( .ip(n4698), .ck(clk), .rb(n12327), .q(
        cache_hit_count[11]) );
  drp_1 \cache_hit_count_reg[10]  ( .ip(n4697), .ck(clk), .rb(n12327), .q(
        cache_hit_count[10]) );
  drp_1 \cache_hit_count_reg[9]  ( .ip(n4696), .ck(clk), .rb(n12327), .q(
        cache_hit_count[9]) );
  drp_1 \cache_hit_count_reg[8]  ( .ip(n4695), .ck(clk), .rb(n12327), .q(
        cache_hit_count[8]) );
  drp_1 \cache_hit_count_reg[7]  ( .ip(n4694), .ck(clk), .rb(n12327), .q(
        cache_hit_count[7]) );
  drp_1 \cache_hit_count_reg[6]  ( .ip(n4693), .ck(clk), .rb(n12327), .q(
        cache_hit_count[6]) );
  drp_1 \cache_hit_count_reg[5]  ( .ip(n4692), .ck(clk), .rb(n12327), .q(
        cache_hit_count[5]) );
  drp_1 \cache_hit_count_reg[4]  ( .ip(n4691), .ck(clk), .rb(n12327), .q(
        cache_hit_count[4]) );
  drp_1 \cache_hit_count_reg[3]  ( .ip(n4690), .ck(clk), .rb(n12327), .q(
        cache_hit_count[3]) );
  drp_1 \cache_hit_count_reg[2]  ( .ip(n4689), .ck(clk), .rb(n12327), .q(
        cache_hit_count[2]) );
  drp_1 \cache_hit_count_reg[1]  ( .ip(n4688), .ck(clk), .rb(n12327), .q(
        cache_hit_count[1]) );
  drp_1 \cache_hit_count_reg[0]  ( .ip(n4687), .ck(clk), .rb(n12327), .q(
        cache_hit_count[0]) );
  invzp_1 \data_rd_tri[4]  ( .ip(n55), .c(N3508), .op(data_rd[4]) );
  invzp_1 \data_rd_tri[5]  ( .ip(n53), .c(N3505), .op(data_rd[5]) );
  invzp_1 \data_rd_tri[8]  ( .ip(n47), .c(N3496), .op(data_rd[8]) );
  invzp_1 \data_rd_tri[10]  ( .ip(n43), .c(N3490), .op(data_rd[10]) );
  invzp_1 \data_rd_tri[12]  ( .ip(n39), .c(N3484), .op(data_rd[12]) );
  invzp_1 \data_rd_tri[17]  ( .ip(n29), .c(N3469), .op(data_rd[17]) );
  invzp_1 \data_rd_tri[19]  ( .ip(n25), .c(N3463), .op(data_rd[19]) );
  invzp_1 \data_rd_tri[20]  ( .ip(n23), .c(N3460), .op(data_rd[20]) );
  invzp_1 \data_rd_tri[22]  ( .ip(n19), .c(N3454), .op(data_rd[22]) );
  invzp_1 \data_rd_tri[25]  ( .ip(n13), .c(N3445), .op(data_rd[25]) );
  invzp_1 \data_rd_tri[26]  ( .ip(n11), .c(N3442), .op(data_rd[26]) );
  invzp_1 \data_rd_tri[27]  ( .ip(n9), .c(N3439), .op(data_rd[27]) );
  invzp_1 \data_rd_tri[28]  ( .ip(n7), .c(N3436), .op(data_rd[28]) );
  invzp_1 \data_rd_tri[30]  ( .ip(n3), .c(N3430), .op(data_rd[30]) );
  invzp_1 \data_rd_tri[31]  ( .ip(n1), .c(N3427), .op(data_rd[31]) );
  invzp_1 \data_rd_tri[0]  ( .ip(n63), .c(N3520), .op(data_rd[0]) );
  invzp_1 \data_rd_tri[1]  ( .ip(n61), .c(N3517), .op(data_rd[1]) );
  invzp_1 \data_rd_tri[2]  ( .ip(n59), .c(N3514), .op(data_rd[2]) );
  invzp_1 \data_rd_tri[3]  ( .ip(n57), .c(N3511), .op(data_rd[3]) );
  invzp_1 \data_rd_tri[6]  ( .ip(n51), .c(N3502), .op(data_rd[6]) );
  invzp_1 \data_rd_tri[7]  ( .ip(n49), .c(N3499), .op(data_rd[7]) );
  invzp_1 \data_rd_tri[9]  ( .ip(n45), .c(N3493), .op(data_rd[9]) );
  invzp_1 \data_rd_tri[11]  ( .ip(n41), .c(N3487), .op(data_rd[11]) );
  invzp_1 \data_rd_tri[13]  ( .ip(n37), .c(N3481), .op(data_rd[13]) );
  invzp_1 \data_rd_tri[14]  ( .ip(n35), .c(N3478), .op(data_rd[14]) );
  invzp_1 \data_rd_tri[15]  ( .ip(n33), .c(N3475), .op(data_rd[15]) );
  invzp_1 \data_rd_tri[16]  ( .ip(n31), .c(N3472), .op(data_rd[16]) );
  invzp_1 \data_rd_tri[18]  ( .ip(n27), .c(N3466), .op(data_rd[18]) );
  invzp_1 \data_rd_tri[21]  ( .ip(n21), .c(N3457), .op(data_rd[21]) );
  invzp_1 \data_rd_tri[23]  ( .ip(n17), .c(N3451), .op(data_rd[23]) );
  invzp_1 \data_rd_tri[24]  ( .ip(n15), .c(N3448), .op(data_rd[24]) );
  invzp_1 \data_rd_tri[29]  ( .ip(n5), .c(N3433), .op(data_rd[29]) );
  invzp_1 \addr_resp_tri[0]  ( .ip(n127), .c(N3616), .op(addr_resp[0]) );
  invzp_1 \addr_resp_tri[1]  ( .ip(n125), .c(N3613), .op(addr_resp[1]) );
  invzp_1 \addr_resp_tri[8]  ( .ip(n111), .c(N3592), .op(addr_resp[8]) );
  invzp_1 \addr_resp_tri[9]  ( .ip(n109), .c(N3589), .op(addr_resp[9]) );
  invzp_1 \addr_resp_tri[10]  ( .ip(n107), .c(N3586), .op(addr_resp[10]) );
  invzp_1 \addr_resp_tri[11]  ( .ip(n105), .c(N3583), .op(addr_resp[11]) );
  invzp_1 \addr_resp_tri[12]  ( .ip(n103), .c(N3580), .op(addr_resp[12]) );
  invzp_1 \addr_resp_tri[13]  ( .ip(n101), .c(N3577), .op(addr_resp[13]) );
  invzp_1 \addr_resp_tri[14]  ( .ip(n99), .c(N3574), .op(addr_resp[14]) );
  invzp_1 \addr_resp_tri[15]  ( .ip(n97), .c(N3571), .op(addr_resp[15]) );
  invzp_1 \addr_resp_tri[16]  ( .ip(n95), .c(N3568), .op(addr_resp[16]) );
  invzp_1 \addr_resp_tri[17]  ( .ip(n93), .c(N3565), .op(addr_resp[17]) );
  invzp_1 \addr_resp_tri[18]  ( .ip(n91), .c(N3562), .op(addr_resp[18]) );
  invzp_1 \addr_resp_tri[19]  ( .ip(n89), .c(N3559), .op(addr_resp[19]) );
  invzp_1 \addr_resp_tri[20]  ( .ip(n87), .c(N3556), .op(addr_resp[20]) );
  invzp_1 \addr_resp_tri[21]  ( .ip(n85), .c(N3553), .op(addr_resp[21]) );
  invzp_1 \addr_resp_tri[22]  ( .ip(n83), .c(N3550), .op(addr_resp[22]) );
  invzp_1 \addr_resp_tri[23]  ( .ip(n81), .c(N3547), .op(addr_resp[23]) );
  invzp_1 \addr_resp_tri[24]  ( .ip(n79), .c(N3544), .op(addr_resp[24]) );
  invzp_1 \addr_resp_tri[25]  ( .ip(n77), .c(N3541), .op(addr_resp[25]) );
  invzp_1 \addr_resp_tri[26]  ( .ip(n75), .c(N3538), .op(addr_resp[26]) );
  invzp_1 \addr_resp_tri[27]  ( .ip(n73), .c(N3535), .op(addr_resp[27]) );
  invzp_1 \addr_resp_tri[28]  ( .ip(n71), .c(N3532), .op(addr_resp[28]) );
  invzp_1 \addr_resp_tri[29]  ( .ip(n69), .c(N3529), .op(addr_resp[29]) );
  invzp_1 \addr_resp_tri[30]  ( .ip(n67), .c(N3526), .op(addr_resp[30]) );
  invzp_1 \addr_resp_tri[31]  ( .ip(n65), .c(N3523), .op(addr_resp[31]) );
  invzp_1 \addr_resp_tri[2]  ( .ip(n123), .c(N3610), .op(addr_resp[2]) );
  invzp_1 \addr_resp_tri[3]  ( .ip(n121), .c(N3607), .op(addr_resp[3]) );
  invzp_1 \addr_resp_tri[5]  ( .ip(n117), .c(N3601), .op(addr_resp[5]) );
  invzp_1 \addr_resp_tri[4]  ( .ip(n119), .c(N3604), .op(addr_resp[4]) );
  invzp_1 \addr_resp_tri[7]  ( .ip(n113), .c(N3595), .op(addr_resp[7]) );
  invzp_1 \addr_resp_tri[6]  ( .ip(n115), .c(N3598), .op(addr_resp[6]) );
  buf_1 U7396 ( .ip(rst), .op(n12324) );
  inv_1 U7397 ( .ip(n12324), .op(n12322) );
  buf_1 U7398 ( .ip(n12322), .op(n12326) );
  buf_1 U7399 ( .ip(rst), .op(n12334) );
  buf_1 U7400 ( .ip(rst), .op(n12335) );
  buf_1 U7401 ( .ip(rst), .op(n12336) );
  inv_1 U7402 ( .ip(state[3]), .op(n8118) );
  inv_1 U7403 ( .ip(state[2]), .op(n8116) );
  nor2_1 U7404 ( .ip1(state[4]), .ip2(state[0]), .op(n8115) );
  nand4_1 U7405 ( .ip1(n8118), .ip2(n8116), .ip3(n8115), .ip4(state[1]), .op(
        n8131) );
  inv_1 U7406 ( .ip(n8131), .op(n12287) );
  nand2_1 U7407 ( .ip1(n12287), .ip2(hit), .op(n7450) );
  inv_1 U7408 ( .ip(cache_hit_count[0]), .op(n7451) );
  nor2_1 U7409 ( .ip1(n7450), .ip2(n7451), .op(n12320) );
  or2_1 U7410 ( .ip1(n7450), .ip2(n12320), .op(n7453) );
  or2_1 U7411 ( .ip1(n7451), .ip2(n12320), .op(n7452) );
  nand2_1 U7412 ( .ip1(n7453), .ip2(n7452), .op(n4687) );
  nand2_1 U7413 ( .ip1(n12320), .ip2(cache_hit_count[1]), .op(n7454) );
  inv_1 U7414 ( .ip(cache_hit_count[2]), .op(n7455) );
  nor2_1 U7415 ( .ip1(n7454), .ip2(n7455), .op(n12319) );
  or2_1 U7416 ( .ip1(n7454), .ip2(n12319), .op(n7457) );
  or2_1 U7417 ( .ip1(n7455), .ip2(n12319), .op(n7456) );
  nand2_1 U7418 ( .ip1(n7457), .ip2(n7456), .op(n4689) );
  nand2_1 U7419 ( .ip1(n12319), .ip2(cache_hit_count[3]), .op(n7458) );
  inv_1 U7420 ( .ip(cache_hit_count[4]), .op(n7459) );
  nor2_1 U7421 ( .ip1(n7458), .ip2(n7459), .op(n12318) );
  or2_1 U7422 ( .ip1(n7458), .ip2(n12318), .op(n7461) );
  or2_1 U7423 ( .ip1(n7459), .ip2(n12318), .op(n7460) );
  nand2_1 U7424 ( .ip1(n7461), .ip2(n7460), .op(n4691) );
  nand2_1 U7425 ( .ip1(n12318), .ip2(cache_hit_count[5]), .op(n7462) );
  inv_1 U7426 ( .ip(cache_hit_count[6]), .op(n7463) );
  nor2_1 U7427 ( .ip1(n7462), .ip2(n7463), .op(n12317) );
  or2_1 U7428 ( .ip1(n7462), .ip2(n12317), .op(n7465) );
  or2_1 U7429 ( .ip1(n7463), .ip2(n12317), .op(n7464) );
  nand2_1 U7430 ( .ip1(n7465), .ip2(n7464), .op(n4693) );
  inv_1 U7431 ( .ip(cache_hit_count[8]), .op(n7466) );
  and3_1 U7432 ( .ip1(n12317), .ip2(cache_hit_count[7]), .ip3(
        cache_hit_count[8]), .op(n12314) );
  or2_1 U7433 ( .ip1(n7466), .ip2(n12314), .op(n7469) );
  nand2_1 U7434 ( .ip1(n12317), .ip2(cache_hit_count[7]), .op(n7467) );
  or2_1 U7435 ( .ip1(n7467), .ip2(n12314), .op(n7468) );
  nand2_1 U7436 ( .ip1(n7469), .ip2(n7468), .op(n4695) );
  inv_1 U7437 ( .ip(cache_hit_count[10]), .op(n7473) );
  nand2_1 U7438 ( .ip1(cache_hit_count[9]), .ip2(n12314), .op(n7470) );
  nor2_1 U7439 ( .ip1(n7473), .ip2(n7470), .op(n12312) );
  or2_1 U7440 ( .ip1(n7473), .ip2(n12312), .op(n7472) );
  or2_1 U7441 ( .ip1(n7470), .ip2(n12312), .op(n7471) );
  nand2_1 U7442 ( .ip1(n7472), .ip2(n7471), .op(n4697) );
  inv_1 U7443 ( .ip(cache_hit_count[12]), .op(n7475) );
  inv_1 U7444 ( .ip(cache_hit_count[9]), .op(n12315) );
  inv_1 U7445 ( .ip(cache_hit_count[11]), .op(n12313) );
  nor4_1 U7446 ( .ip1(n12315), .ip2(n7473), .ip3(n12313), .ip4(n7475), .op(
        n7474) );
  nand4_1 U7447 ( .ip1(n12317), .ip2(cache_hit_count[7]), .ip3(
        cache_hit_count[8]), .ip4(n7474), .op(n7480) );
  inv_1 U7448 ( .ip(n7480), .op(n7476) );
  or2_1 U7449 ( .ip1(n7475), .ip2(n7476), .op(n7479) );
  nand2_1 U7450 ( .ip1(cache_hit_count[11]), .ip2(n12312), .op(n7477) );
  or2_1 U7451 ( .ip1(n7477), .ip2(n7476), .op(n7478) );
  nand2_1 U7452 ( .ip1(n7479), .ip2(n7478), .op(n4699) );
  inv_1 U7453 ( .ip(cache_hit_count[13]), .op(n7481) );
  nor2_1 U7454 ( .ip1(n7480), .ip2(n7481), .op(n12311) );
  or2_1 U7455 ( .ip1(n7480), .ip2(n12311), .op(n7483) );
  or2_1 U7456 ( .ip1(n7481), .ip2(n12311), .op(n7482) );
  nand2_1 U7457 ( .ip1(n7483), .ip2(n7482), .op(n4700) );
  nand2_1 U7458 ( .ip1(n12311), .ip2(cache_hit_count[14]), .op(n7484) );
  inv_1 U7459 ( .ip(cache_hit_count[15]), .op(n7485) );
  nor2_1 U7460 ( .ip1(n7484), .ip2(n7485), .op(n12308) );
  or2_1 U7461 ( .ip1(n7484), .ip2(n12308), .op(n7487) );
  or2_1 U7462 ( .ip1(n7485), .ip2(n12308), .op(n7486) );
  nand2_1 U7463 ( .ip1(n7487), .ip2(n7486), .op(n4702) );
  nand2_1 U7464 ( .ip1(n12308), .ip2(cache_hit_count[16]), .op(n12307) );
  inv_1 U7465 ( .ip(cache_hit_count[17]), .op(n7488) );
  nor2_1 U7466 ( .ip1(n12307), .ip2(n7488), .op(n12305) );
  or2_1 U7467 ( .ip1(n12307), .ip2(n12305), .op(n7490) );
  or2_1 U7468 ( .ip1(n7488), .ip2(n12305), .op(n7489) );
  nand2_1 U7469 ( .ip1(n7490), .ip2(n7489), .op(n4704) );
  inv_1 U7470 ( .ip(cache_hit_count[19]), .op(n7491) );
  nand2_1 U7471 ( .ip1(cache_hit_count[18]), .ip2(n12305), .op(n12298) );
  nor2_1 U7472 ( .ip1(n7491), .ip2(n12298), .op(n12302) );
  or2_1 U7473 ( .ip1(n7491), .ip2(n12302), .op(n7493) );
  or2_1 U7474 ( .ip1(n12298), .ip2(n12302), .op(n7492) );
  nand2_1 U7475 ( .ip1(n7493), .ip2(n7492), .op(n4706) );
  nand2_1 U7476 ( .ip1(cache_hit_count[19]), .ip2(cache_hit_count[20]), .op(
        n12299) );
  nor2_1 U7477 ( .ip1(n12307), .ip2(n12299), .op(n7494) );
  nand4_1 U7478 ( .ip1(cache_hit_count[21]), .ip2(cache_hit_count[17]), .ip3(
        cache_hit_count[18]), .ip4(n7494), .op(n12297) );
  inv_1 U7479 ( .ip(cache_hit_count[22]), .op(n7495) );
  nor2_1 U7480 ( .ip1(n12297), .ip2(n7495), .op(n12296) );
  or2_1 U7481 ( .ip1(n12297), .ip2(n12296), .op(n7497) );
  or2_1 U7482 ( .ip1(n7495), .ip2(n12296), .op(n7496) );
  nand2_1 U7483 ( .ip1(n7497), .ip2(n7496), .op(n4709) );
  nand2_1 U7484 ( .ip1(n12296), .ip2(cache_hit_count[23]), .op(n7498) );
  inv_1 U7485 ( .ip(cache_hit_count[24]), .op(n7499) );
  nor2_1 U7486 ( .ip1(n7498), .ip2(n7499), .op(n12295) );
  or2_1 U7487 ( .ip1(n7498), .ip2(n12295), .op(n7501) );
  or2_1 U7488 ( .ip1(n7499), .ip2(n12295), .op(n7500) );
  nand2_1 U7489 ( .ip1(n7501), .ip2(n7500), .op(n4711) );
  nand2_1 U7490 ( .ip1(n12295), .ip2(cache_hit_count[25]), .op(n7502) );
  inv_1 U7491 ( .ip(cache_hit_count[26]), .op(n7503) );
  nor2_1 U7492 ( .ip1(n7502), .ip2(n7503), .op(n12294) );
  or2_1 U7493 ( .ip1(n7502), .ip2(n12294), .op(n7505) );
  or2_1 U7494 ( .ip1(n7503), .ip2(n12294), .op(n7504) );
  nand2_1 U7495 ( .ip1(n7505), .ip2(n7504), .op(n4713) );
  nand2_1 U7496 ( .ip1(n12294), .ip2(cache_hit_count[27]), .op(n7506) );
  inv_1 U7497 ( .ip(cache_hit_count[28]), .op(n7507) );
  nor2_1 U7498 ( .ip1(n7506), .ip2(n7507), .op(n12293) );
  or2_1 U7499 ( .ip1(n7506), .ip2(n12293), .op(n7509) );
  or2_1 U7500 ( .ip1(n7507), .ip2(n12293), .op(n7508) );
  nand2_1 U7501 ( .ip1(n7509), .ip2(n7508), .op(n4715) );
  nand3_1 U7502 ( .ip1(n12287), .ip2(miss), .ip3(cache_miss_count[0]), .op(
        n7510) );
  inv_1 U7503 ( .ip(cache_miss_count[1]), .op(n7511) );
  nor2_1 U7504 ( .ip1(n7510), .ip2(n7511), .op(n12286) );
  or2_1 U7505 ( .ip1(n7510), .ip2(n12286), .op(n7513) );
  or2_1 U7506 ( .ip1(n7511), .ip2(n12286), .op(n7512) );
  nand2_1 U7507 ( .ip1(n7513), .ip2(n7512), .op(n4720) );
  nand2_1 U7508 ( .ip1(n12286), .ip2(cache_miss_count[2]), .op(n7514) );
  inv_1 U7509 ( .ip(cache_miss_count[3]), .op(n7515) );
  nor2_1 U7510 ( .ip1(n7514), .ip2(n7515), .op(n12285) );
  or2_1 U7511 ( .ip1(n7514), .ip2(n12285), .op(n7517) );
  or2_1 U7512 ( .ip1(n7515), .ip2(n12285), .op(n7516) );
  nand2_1 U7513 ( .ip1(n7517), .ip2(n7516), .op(n4722) );
  nand2_1 U7514 ( .ip1(n12285), .ip2(cache_miss_count[4]), .op(n7518) );
  inv_1 U7515 ( .ip(cache_miss_count[5]), .op(n7519) );
  nor2_1 U7516 ( .ip1(n7518), .ip2(n7519), .op(n12282) );
  or2_1 U7517 ( .ip1(n7518), .ip2(n12282), .op(n7521) );
  or2_1 U7518 ( .ip1(n7519), .ip2(n12282), .op(n7520) );
  nand2_1 U7519 ( .ip1(n7521), .ip2(n7520), .op(n4724) );
  nand2_1 U7520 ( .ip1(n12282), .ip2(cache_miss_count[6]), .op(n12281) );
  inv_1 U7521 ( .ip(cache_miss_count[7]), .op(n7522) );
  nor2_1 U7522 ( .ip1(n12281), .ip2(n7522), .op(n12279) );
  or2_1 U7523 ( .ip1(n12281), .ip2(n12279), .op(n7524) );
  or2_1 U7524 ( .ip1(n7522), .ip2(n12279), .op(n7523) );
  nand2_1 U7525 ( .ip1(n7524), .ip2(n7523), .op(n4726) );
  inv_1 U7526 ( .ip(cache_miss_count[9]), .op(n7525) );
  nand2_1 U7527 ( .ip1(cache_miss_count[8]), .ip2(n12279), .op(n7526) );
  nor2_1 U7528 ( .ip1(n7525), .ip2(n7526), .op(n12277) );
  or2_1 U7529 ( .ip1(n7525), .ip2(n12277), .op(n7528) );
  or2_1 U7530 ( .ip1(n7526), .ip2(n12277), .op(n7527) );
  nand2_1 U7531 ( .ip1(n7528), .ip2(n7527), .op(n4728) );
  inv_1 U7532 ( .ip(cache_miss_count[11]), .op(n7529) );
  nand2_1 U7533 ( .ip1(cache_miss_count[10]), .ip2(n12277), .op(n7530) );
  nor2_1 U7534 ( .ip1(n7529), .ip2(n7530), .op(n12275) );
  or2_1 U7535 ( .ip1(n7529), .ip2(n12275), .op(n7532) );
  or2_1 U7536 ( .ip1(n7530), .ip2(n12275), .op(n7531) );
  nand2_1 U7537 ( .ip1(n7532), .ip2(n7531), .op(n4730) );
  inv_1 U7538 ( .ip(cache_miss_count[13]), .op(n7533) );
  nand2_1 U7539 ( .ip1(cache_miss_count[12]), .ip2(n12275), .op(n7534) );
  nor2_1 U7540 ( .ip1(n7533), .ip2(n7534), .op(n12273) );
  or2_1 U7541 ( .ip1(n7533), .ip2(n12273), .op(n7536) );
  or2_1 U7542 ( .ip1(n7534), .ip2(n12273), .op(n7535) );
  nand2_1 U7543 ( .ip1(n7536), .ip2(n7535), .op(n4732) );
  inv_1 U7544 ( .ip(cache_miss_count[15]), .op(n7537) );
  nand2_1 U7545 ( .ip1(cache_miss_count[14]), .ip2(n12273), .op(n7538) );
  nor2_1 U7546 ( .ip1(n7537), .ip2(n7538), .op(n12270) );
  or2_1 U7547 ( .ip1(n7537), .ip2(n12270), .op(n7540) );
  or2_1 U7548 ( .ip1(n7538), .ip2(n12270), .op(n7539) );
  nand2_1 U7549 ( .ip1(n7540), .ip2(n7539), .op(n4734) );
  nand4_1 U7550 ( .ip1(cache_miss_count[7]), .ip2(cache_miss_count[8]), .ip3(
        cache_miss_count[9]), .ip4(cache_miss_count[10]), .op(n7543) );
  nand4_1 U7551 ( .ip1(cache_miss_count[11]), .ip2(cache_miss_count[12]), 
        .ip3(cache_miss_count[13]), .ip4(cache_miss_count[14]), .op(n7542) );
  nand4_1 U7552 ( .ip1(cache_miss_count[15]), .ip2(cache_miss_count[16]), 
        .ip3(cache_miss_count[17]), .ip4(cache_miss_count[18]), .op(n7541) );
  nor4_1 U7553 ( .ip1(n12281), .ip2(n7543), .ip3(n7542), .ip4(n7541), .op(
        n12266) );
  nand2_1 U7554 ( .ip1(n12266), .ip2(cache_miss_count[19]), .op(n7544) );
  inv_1 U7555 ( .ip(cache_miss_count[20]), .op(n7545) );
  nor2_1 U7556 ( .ip1(n7544), .ip2(n7545), .op(n12265) );
  or2_1 U7557 ( .ip1(n7544), .ip2(n12265), .op(n7547) );
  or2_1 U7558 ( .ip1(n7545), .ip2(n12265), .op(n7546) );
  nand2_1 U7559 ( .ip1(n7547), .ip2(n7546), .op(n4739) );
  nand2_1 U7560 ( .ip1(n12265), .ip2(cache_miss_count[21]), .op(n7548) );
  inv_1 U7561 ( .ip(cache_miss_count[22]), .op(n7549) );
  nor2_1 U7562 ( .ip1(n7548), .ip2(n7549), .op(n12264) );
  or2_1 U7563 ( .ip1(n7548), .ip2(n12264), .op(n7551) );
  or2_1 U7564 ( .ip1(n7549), .ip2(n12264), .op(n7550) );
  nand2_1 U7565 ( .ip1(n7551), .ip2(n7550), .op(n4741) );
  nand2_1 U7566 ( .ip1(n12264), .ip2(cache_miss_count[23]), .op(n7552) );
  inv_1 U7567 ( .ip(cache_miss_count[24]), .op(n7553) );
  nor2_1 U7568 ( .ip1(n7552), .ip2(n7553), .op(n12263) );
  or2_1 U7569 ( .ip1(n7552), .ip2(n12263), .op(n7555) );
  or2_1 U7570 ( .ip1(n7553), .ip2(n12263), .op(n7554) );
  nand2_1 U7571 ( .ip1(n7555), .ip2(n7554), .op(n4743) );
  nand2_1 U7572 ( .ip1(n12263), .ip2(cache_miss_count[25]), .op(n7556) );
  inv_1 U7573 ( .ip(cache_miss_count[26]), .op(n7557) );
  nor2_1 U7574 ( .ip1(n7556), .ip2(n7557), .op(n12262) );
  or2_1 U7575 ( .ip1(n7556), .ip2(n12262), .op(n7559) );
  or2_1 U7576 ( .ip1(n7557), .ip2(n12262), .op(n7558) );
  nand2_1 U7577 ( .ip1(n7559), .ip2(n7558), .op(n4745) );
  nand2_1 U7578 ( .ip1(n12262), .ip2(cache_miss_count[27]), .op(n7560) );
  inv_1 U7579 ( .ip(cache_miss_count[28]), .op(n7561) );
  nor2_1 U7580 ( .ip1(n7560), .ip2(n7561), .op(n12261) );
  or2_1 U7581 ( .ip1(n7560), .ip2(n12261), .op(n7563) );
  or2_1 U7582 ( .ip1(n7561), .ip2(n12261), .op(n7562) );
  nand2_1 U7583 ( .ip1(n7563), .ip2(n7562), .op(n4747) );
  inv_1 U7584 ( .ip(mem_data_cnt[3]), .op(n11438) );
  inv_1 U7585 ( .ip(mem_data_cnt[2]), .op(n11433) );
  nor2_1 U7586 ( .ip1(n11438), .ip2(n11433), .op(N3698) );
  nor2_1 U7587 ( .ip1(wr), .ip2(rd), .op(n7727) );
  inv_1 U7588 ( .ip(state[0]), .op(n7564) );
  nor4_1 U7589 ( .ip1(state[4]), .ip2(state[1]), .ip3(n7727), .ip4(n7564), 
        .op(n7565) );
  nand3_1 U7590 ( .ip1(n7565), .ip2(n8118), .ip3(n8116), .op(n8130) );
  inv_1 U7591 ( .ip(miss), .op(n8119) );
  inv_1 U7592 ( .ip(hit), .op(n11357) );
  nand4_1 U7593 ( .ip1(n12287), .ip2(valid), .ip3(n8119), .ip4(n11357), .op(
        n7566) );
  nand2_1 U7594 ( .ip1(n8130), .ip2(n7566), .op(next_state[1]) );
  nand2_1 U7595 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .op(n7584) );
  nor3_1 U7596 ( .ip1(addr_req[7]), .ip2(addr_req[6]), .ip3(n7584), .op(n10931) );
  nand2_1 U7597 ( .ip1(\cache_tag[3][14] ), .ip2(n10931), .op(n7570) );
  inv_1 U7598 ( .ip(addr_req[6]), .op(n7576) );
  or2_1 U7599 ( .ip1(n7576), .ip2(addr_req[7]), .op(n7577) );
  nor3_1 U7600 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .ip3(n7577), .op(n10948) );
  nand2_1 U7601 ( .ip1(\cache_tag[4][14] ), .ip2(n10948), .op(n7569) );
  nor2_1 U7602 ( .ip1(n7584), .ip2(n7577), .op(n10933) );
  nand2_1 U7603 ( .ip1(\cache_tag[7][14] ), .ip2(n10933), .op(n7568) );
  inv_1 U7604 ( .ip(addr_req[4]), .op(n7571) );
  or2_1 U7605 ( .ip1(n7571), .ip2(addr_req[5]), .op(n7586) );
  nand2_1 U7606 ( .ip1(addr_req[7]), .ip2(addr_req[6]), .op(n7583) );
  nor2_1 U7607 ( .ip1(n7586), .ip2(n7583), .op(n10949) );
  nand2_1 U7608 ( .ip1(\cache_tag[13][14] ), .ip2(n10949), .op(n7567) );
  nand4_1 U7609 ( .ip1(n7570), .ip2(n7569), .ip3(n7568), .ip4(n7567), .op(
        n7594) );
  nand2_1 U7610 ( .ip1(addr_req[5]), .ip2(n7571), .op(n7578) );
  nor2_1 U7611 ( .ip1(n7583), .ip2(n7578), .op(n10938) );
  nand2_1 U7612 ( .ip1(\cache_tag[14][14] ), .ip2(n10938), .op(n7575) );
  nor3_1 U7613 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .ip3(n7583), .op(n10939) );
  nand2_1 U7614 ( .ip1(\cache_tag[12][14] ), .ip2(n10939), .op(n7574) );
  nor3_1 U7615 ( .ip1(addr_req[7]), .ip2(addr_req[6]), .ip3(n7578), .op(n10925) );
  nand2_1 U7616 ( .ip1(\cache_tag[2][14] ), .ip2(n10925), .op(n7573) );
  nor4_1 U7617 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .ip3(addr_req[7]), 
        .ip4(addr_req[6]), .op(n10946) );
  nand2_1 U7618 ( .ip1(\cache_tag[0][14] ), .ip2(n10946), .op(n7572) );
  nand4_1 U7619 ( .ip1(n7575), .ip2(n7574), .ip3(n7573), .ip4(n7572), .op(
        n7593) );
  nor2_1 U7620 ( .ip1(n7577), .ip2(n7578), .op(n10924) );
  nand2_1 U7621 ( .ip1(\cache_tag[6][14] ), .ip2(n10924), .op(n7582) );
  nand2_1 U7622 ( .ip1(addr_req[7]), .ip2(n7576), .op(n7585) );
  nor2_1 U7623 ( .ip1(n7584), .ip2(n7585), .op(n10941) );
  nand2_1 U7624 ( .ip1(\cache_tag[11][14] ), .ip2(n10941), .op(n7581) );
  nor2_1 U7625 ( .ip1(n7577), .ip2(n7586), .op(n10947) );
  nand2_1 U7626 ( .ip1(\cache_tag[5][14] ), .ip2(n10947), .op(n7580) );
  nor2_1 U7627 ( .ip1(n7578), .ip2(n7585), .op(n10922) );
  nand2_1 U7628 ( .ip1(\cache_tag[10][14] ), .ip2(n10922), .op(n7579) );
  nand4_1 U7629 ( .ip1(n7582), .ip2(n7581), .ip3(n7580), .ip4(n7579), .op(
        n7592) );
  nor2_1 U7630 ( .ip1(n7584), .ip2(n7583), .op(n10940) );
  nand2_1 U7631 ( .ip1(\cache_tag[15][14] ), .ip2(n10940), .op(n7590) );
  nor2_1 U7632 ( .ip1(n7586), .ip2(n7585), .op(n10923) );
  nand2_1 U7633 ( .ip1(\cache_tag[9][14] ), .ip2(n10923), .op(n7589) );
  nor3_1 U7634 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .ip3(n7585), .op(n10932) );
  nand2_1 U7635 ( .ip1(\cache_tag[8][14] ), .ip2(n10932), .op(n7588) );
  nor3_1 U7636 ( .ip1(addr_req[7]), .ip2(addr_req[6]), .ip3(n7586), .op(n10930) );
  nand2_1 U7637 ( .ip1(\cache_tag[1][14] ), .ip2(n10930), .op(n7587) );
  nand4_1 U7638 ( .ip1(n7590), .ip2(n7589), .ip3(n7588), .ip4(n7587), .op(
        n7591) );
  nor4_1 U7639 ( .ip1(n7594), .ip2(n7593), .ip3(n7592), .ip4(n7591), .op(n7595) );
  xor2_1 U7640 ( .ip1(addr_req[22]), .ip2(n7595), .op(n7662) );
  nand2_1 U7641 ( .ip1(n10933), .ip2(\cache_tag[7][9] ), .op(n7599) );
  nand2_1 U7642 ( .ip1(n10941), .ip2(\cache_tag[11][9] ), .op(n7598) );
  nand2_1 U7643 ( .ip1(n10940), .ip2(\cache_tag[15][9] ), .op(n7597) );
  nand2_1 U7644 ( .ip1(n10948), .ip2(\cache_tag[4][9] ), .op(n7596) );
  nand4_1 U7645 ( .ip1(n7599), .ip2(n7598), .ip3(n7597), .ip4(n7596), .op(
        n7615) );
  nand2_1 U7646 ( .ip1(n10924), .ip2(\cache_tag[6][9] ), .op(n7603) );
  nand2_1 U7647 ( .ip1(n10930), .ip2(\cache_tag[1][9] ), .op(n7602) );
  nand2_1 U7648 ( .ip1(n10949), .ip2(\cache_tag[13][9] ), .op(n7601) );
  nand2_1 U7649 ( .ip1(n10922), .ip2(\cache_tag[10][9] ), .op(n7600) );
  nand4_1 U7650 ( .ip1(n7603), .ip2(n7602), .ip3(n7601), .ip4(n7600), .op(
        n7614) );
  nand2_1 U7651 ( .ip1(n10931), .ip2(\cache_tag[3][9] ), .op(n7607) );
  nand2_1 U7652 ( .ip1(n10938), .ip2(\cache_tag[14][9] ), .op(n7606) );
  nand2_1 U7653 ( .ip1(n10946), .ip2(\cache_tag[0][9] ), .op(n7605) );
  nand2_1 U7654 ( .ip1(n10939), .ip2(\cache_tag[12][9] ), .op(n7604) );
  nand4_1 U7655 ( .ip1(n7607), .ip2(n7606), .ip3(n7605), .ip4(n7604), .op(
        n7613) );
  nand2_1 U7656 ( .ip1(n10923), .ip2(\cache_tag[9][9] ), .op(n7611) );
  nand2_1 U7657 ( .ip1(n10947), .ip2(\cache_tag[5][9] ), .op(n7610) );
  nand2_1 U7658 ( .ip1(n10932), .ip2(\cache_tag[8][9] ), .op(n7609) );
  nand2_1 U7659 ( .ip1(n10925), .ip2(\cache_tag[2][9] ), .op(n7608) );
  nand4_1 U7660 ( .ip1(n7611), .ip2(n7610), .ip3(n7609), .ip4(n7608), .op(
        n7612) );
  nor4_1 U7661 ( .ip1(n7615), .ip2(n7614), .ip3(n7613), .ip4(n7612), .op(n7616) );
  xor2_1 U7662 ( .ip1(addr_req[17]), .ip2(n7616), .op(n7661) );
  nand2_1 U7663 ( .ip1(n10924), .ip2(\cache_tag[6][13] ), .op(n7620) );
  nand2_1 U7664 ( .ip1(n10933), .ip2(\cache_tag[7][13] ), .op(n7619) );
  nand2_1 U7665 ( .ip1(n10922), .ip2(\cache_tag[10][13] ), .op(n7618) );
  nand2_1 U7666 ( .ip1(n10940), .ip2(\cache_tag[15][13] ), .op(n7617) );
  nand4_1 U7667 ( .ip1(n7620), .ip2(n7619), .ip3(n7618), .ip4(n7617), .op(
        n7636) );
  nand2_1 U7668 ( .ip1(n10939), .ip2(\cache_tag[12][13] ), .op(n7624) );
  nand2_1 U7669 ( .ip1(n10923), .ip2(\cache_tag[9][13] ), .op(n7623) );
  nand2_1 U7670 ( .ip1(n10930), .ip2(\cache_tag[1][13] ), .op(n7622) );
  nand2_1 U7671 ( .ip1(n10949), .ip2(\cache_tag[13][13] ), .op(n7621) );
  nand4_1 U7672 ( .ip1(n7624), .ip2(n7623), .ip3(n7622), .ip4(n7621), .op(
        n7635) );
  nand2_1 U7673 ( .ip1(n10925), .ip2(\cache_tag[2][13] ), .op(n7628) );
  nand2_1 U7674 ( .ip1(n10938), .ip2(\cache_tag[14][13] ), .op(n7627) );
  nand2_1 U7675 ( .ip1(n10948), .ip2(\cache_tag[4][13] ), .op(n7626) );
  nand2_1 U7676 ( .ip1(n10931), .ip2(\cache_tag[3][13] ), .op(n7625) );
  nand4_1 U7677 ( .ip1(n7628), .ip2(n7627), .ip3(n7626), .ip4(n7625), .op(
        n7634) );
  nand2_1 U7678 ( .ip1(n10941), .ip2(\cache_tag[11][13] ), .op(n7632) );
  nand2_1 U7679 ( .ip1(n10946), .ip2(\cache_tag[0][13] ), .op(n7631) );
  nand2_1 U7680 ( .ip1(n10932), .ip2(\cache_tag[8][13] ), .op(n7630) );
  nand2_1 U7681 ( .ip1(n10947), .ip2(\cache_tag[5][13] ), .op(n7629) );
  nand4_1 U7682 ( .ip1(n7632), .ip2(n7631), .ip3(n7630), .ip4(n7629), .op(
        n7633) );
  nor4_1 U7683 ( .ip1(n7636), .ip2(n7635), .ip3(n7634), .ip4(n7633), .op(n7637) );
  xor2_1 U7684 ( .ip1(addr_req[21]), .ip2(n7637), .op(n7660) );
  nand2_1 U7685 ( .ip1(n10923), .ip2(\cache_tag[9][20] ), .op(n7641) );
  nand2_1 U7686 ( .ip1(n10932), .ip2(\cache_tag[8][20] ), .op(n7640) );
  nand2_1 U7687 ( .ip1(n10948), .ip2(\cache_tag[4][20] ), .op(n7639) );
  nand2_1 U7688 ( .ip1(n10938), .ip2(\cache_tag[14][20] ), .op(n7638) );
  nand4_1 U7689 ( .ip1(n7641), .ip2(n7640), .ip3(n7639), .ip4(n7638), .op(
        n7657) );
  nand2_1 U7690 ( .ip1(n10940), .ip2(\cache_tag[15][20] ), .op(n7645) );
  nand2_1 U7691 ( .ip1(n10949), .ip2(\cache_tag[13][20] ), .op(n7644) );
  nand2_1 U7692 ( .ip1(n10924), .ip2(\cache_tag[6][20] ), .op(n7643) );
  nand2_1 U7693 ( .ip1(n10947), .ip2(\cache_tag[5][20] ), .op(n7642) );
  nand4_1 U7694 ( .ip1(n7645), .ip2(n7644), .ip3(n7643), .ip4(n7642), .op(
        n7656) );
  nand2_1 U7695 ( .ip1(n10946), .ip2(\cache_tag[0][20] ), .op(n7649) );
  nand2_1 U7696 ( .ip1(n10939), .ip2(\cache_tag[12][20] ), .op(n7648) );
  nand2_1 U7697 ( .ip1(n10931), .ip2(\cache_tag[3][20] ), .op(n7647) );
  nand2_1 U7698 ( .ip1(n10941), .ip2(\cache_tag[11][20] ), .op(n7646) );
  nand4_1 U7699 ( .ip1(n7649), .ip2(n7648), .ip3(n7647), .ip4(n7646), .op(
        n7655) );
  nand2_1 U7700 ( .ip1(n10922), .ip2(\cache_tag[10][20] ), .op(n7653) );
  nand2_1 U7701 ( .ip1(n10925), .ip2(\cache_tag[2][20] ), .op(n7652) );
  nand2_1 U7702 ( .ip1(n10930), .ip2(\cache_tag[1][20] ), .op(n7651) );
  nand2_1 U7703 ( .ip1(n10933), .ip2(\cache_tag[7][20] ), .op(n7650) );
  nand4_1 U7704 ( .ip1(n7653), .ip2(n7652), .ip3(n7651), .ip4(n7650), .op(
        n7654) );
  nor4_1 U7705 ( .ip1(n7657), .ip2(n7656), .ip3(n7655), .ip4(n7654), .op(n7658) );
  xor2_1 U7706 ( .ip1(addr_req[28]), .ip2(n7658), .op(n7659) );
  nand4_1 U7707 ( .ip1(n7662), .ip2(n7661), .ip3(n7660), .ip4(n7659), .op(
        n8112) );
  inv_1 U7708 ( .ip(addr_req[23]), .op(n7684) );
  nand2_1 U7709 ( .ip1(n10941), .ip2(\cache_tag[11][15] ), .op(n7666) );
  nand2_1 U7710 ( .ip1(n10939), .ip2(\cache_tag[12][15] ), .op(n7665) );
  nand2_1 U7711 ( .ip1(n10925), .ip2(\cache_tag[2][15] ), .op(n7664) );
  nand2_1 U7712 ( .ip1(n10930), .ip2(\cache_tag[1][15] ), .op(n7663) );
  nand4_1 U7713 ( .ip1(n7666), .ip2(n7665), .ip3(n7664), .ip4(n7663), .op(
        n7682) );
  nand2_1 U7714 ( .ip1(n10931), .ip2(\cache_tag[3][15] ), .op(n7670) );
  nand2_1 U7715 ( .ip1(n10933), .ip2(\cache_tag[7][15] ), .op(n7669) );
  nand2_1 U7716 ( .ip1(n10940), .ip2(\cache_tag[15][15] ), .op(n7668) );
  nand2_1 U7717 ( .ip1(n10938), .ip2(\cache_tag[14][15] ), .op(n7667) );
  nand4_1 U7718 ( .ip1(n7670), .ip2(n7669), .ip3(n7668), .ip4(n7667), .op(
        n7681) );
  nand2_1 U7719 ( .ip1(n10948), .ip2(\cache_tag[4][15] ), .op(n7674) );
  nand2_1 U7720 ( .ip1(n10947), .ip2(\cache_tag[5][15] ), .op(n7673) );
  nand2_1 U7721 ( .ip1(n10932), .ip2(\cache_tag[8][15] ), .op(n7672) );
  nand2_1 U7722 ( .ip1(n10924), .ip2(\cache_tag[6][15] ), .op(n7671) );
  nand4_1 U7723 ( .ip1(n7674), .ip2(n7673), .ip3(n7672), .ip4(n7671), .op(
        n7680) );
  nand2_1 U7724 ( .ip1(n10949), .ip2(\cache_tag[13][15] ), .op(n7678) );
  nand2_1 U7725 ( .ip1(n10923), .ip2(\cache_tag[9][15] ), .op(n7677) );
  nand2_1 U7726 ( .ip1(n10922), .ip2(\cache_tag[10][15] ), .op(n7676) );
  nand2_1 U7727 ( .ip1(n10946), .ip2(\cache_tag[0][15] ), .op(n7675) );
  nand4_1 U7728 ( .ip1(n7678), .ip2(n7677), .ip3(n7676), .ip4(n7675), .op(
        n7679) );
  nor4_1 U7729 ( .ip1(n7682), .ip2(n7681), .ip3(n7680), .ip4(n7679), .op(n7683) );
  mux2_1 U7730 ( .ip1(n7684), .ip2(addr_req[23]), .s(n7683), .op(n8111) );
  nand2_1 U7731 ( .ip1(n10923), .ip2(\cache_tag[9][12] ), .op(n7688) );
  nand2_1 U7732 ( .ip1(n10939), .ip2(\cache_tag[12][12] ), .op(n7687) );
  nand2_1 U7733 ( .ip1(n10947), .ip2(\cache_tag[5][12] ), .op(n7686) );
  nand2_1 U7734 ( .ip1(n10930), .ip2(\cache_tag[1][12] ), .op(n7685) );
  nand4_1 U7735 ( .ip1(n7688), .ip2(n7687), .ip3(n7686), .ip4(n7685), .op(
        n7704) );
  nand2_1 U7736 ( .ip1(n10924), .ip2(\cache_tag[6][12] ), .op(n7692) );
  nand2_1 U7737 ( .ip1(n10938), .ip2(\cache_tag[14][12] ), .op(n7691) );
  nand2_1 U7738 ( .ip1(n10932), .ip2(\cache_tag[8][12] ), .op(n7690) );
  nand2_1 U7739 ( .ip1(n10925), .ip2(\cache_tag[2][12] ), .op(n7689) );
  nand4_1 U7740 ( .ip1(n7692), .ip2(n7691), .ip3(n7690), .ip4(n7689), .op(
        n7703) );
  nand2_1 U7741 ( .ip1(n10940), .ip2(\cache_tag[15][12] ), .op(n7696) );
  nand2_1 U7742 ( .ip1(n10946), .ip2(\cache_tag[0][12] ), .op(n7695) );
  nand2_1 U7743 ( .ip1(n10949), .ip2(\cache_tag[13][12] ), .op(n7694) );
  nand2_1 U7744 ( .ip1(n10941), .ip2(\cache_tag[11][12] ), .op(n7693) );
  nand4_1 U7745 ( .ip1(n7696), .ip2(n7695), .ip3(n7694), .ip4(n7693), .op(
        n7702) );
  nand2_1 U7746 ( .ip1(n10933), .ip2(\cache_tag[7][12] ), .op(n7700) );
  nand2_1 U7747 ( .ip1(n10948), .ip2(\cache_tag[4][12] ), .op(n7699) );
  nand2_1 U7748 ( .ip1(n10922), .ip2(\cache_tag[10][12] ), .op(n7698) );
  nand2_1 U7749 ( .ip1(n10931), .ip2(\cache_tag[3][12] ), .op(n7697) );
  nand4_1 U7750 ( .ip1(n7700), .ip2(n7699), .ip3(n7698), .ip4(n7697), .op(
        n7701) );
  nor4_1 U7751 ( .ip1(n7704), .ip2(n7703), .ip3(n7702), .ip4(n7701), .op(n7705) );
  xor2_1 U7752 ( .ip1(addr_req[20]), .ip2(n7705), .op(n7752) );
  nand2_1 U7753 ( .ip1(n10939), .ip2(\cache_tag[12][11] ), .op(n7709) );
  nand2_1 U7754 ( .ip1(n10925), .ip2(\cache_tag[2][11] ), .op(n7708) );
  nand2_1 U7755 ( .ip1(n10940), .ip2(\cache_tag[15][11] ), .op(n7707) );
  nand2_1 U7756 ( .ip1(n10948), .ip2(\cache_tag[4][11] ), .op(n7706) );
  nand4_1 U7757 ( .ip1(n7709), .ip2(n7708), .ip3(n7707), .ip4(n7706), .op(
        n7725) );
  nand2_1 U7758 ( .ip1(n10931), .ip2(\cache_tag[3][11] ), .op(n7713) );
  nand2_1 U7759 ( .ip1(n10949), .ip2(\cache_tag[13][11] ), .op(n7712) );
  nand2_1 U7760 ( .ip1(n10932), .ip2(\cache_tag[8][11] ), .op(n7711) );
  nand2_1 U7761 ( .ip1(n10930), .ip2(\cache_tag[1][11] ), .op(n7710) );
  nand4_1 U7762 ( .ip1(n7713), .ip2(n7712), .ip3(n7711), .ip4(n7710), .op(
        n7724) );
  nand2_1 U7763 ( .ip1(n10924), .ip2(\cache_tag[6][11] ), .op(n7717) );
  nand2_1 U7764 ( .ip1(n10922), .ip2(\cache_tag[10][11] ), .op(n7716) );
  nand2_1 U7765 ( .ip1(n10946), .ip2(\cache_tag[0][11] ), .op(n7715) );
  nand2_1 U7766 ( .ip1(n10933), .ip2(\cache_tag[7][11] ), .op(n7714) );
  nand4_1 U7767 ( .ip1(n7717), .ip2(n7716), .ip3(n7715), .ip4(n7714), .op(
        n7723) );
  nand2_1 U7768 ( .ip1(n10923), .ip2(\cache_tag[9][11] ), .op(n7721) );
  nand2_1 U7769 ( .ip1(n10941), .ip2(\cache_tag[11][11] ), .op(n7720) );
  nand2_1 U7770 ( .ip1(n10938), .ip2(\cache_tag[14][11] ), .op(n7719) );
  nand2_1 U7771 ( .ip1(n10947), .ip2(\cache_tag[5][11] ), .op(n7718) );
  nand4_1 U7772 ( .ip1(n7721), .ip2(n7720), .ip3(n7719), .ip4(n7718), .op(
        n7722) );
  nor4_1 U7773 ( .ip1(n7725), .ip2(n7724), .ip3(n7723), .ip4(n7722), .op(n7726) );
  xor2_1 U7774 ( .ip1(addr_req[19]), .ip2(n7726), .op(n7751) );
  inv_1 U7775 ( .ip(next_state[1]), .op(n10900) );
  nor2_1 U7776 ( .ip1(n7727), .ip2(n10900), .op(n7728) );
  inv_1 U7777 ( .ip(n7728), .op(n11361) );
  inv_1 U7778 ( .ip(n11361), .op(n11358) );
  nand2_1 U7779 ( .ip1(n10933), .ip2(\cache_tag[7][18] ), .op(n7732) );
  nand2_1 U7780 ( .ip1(n10947), .ip2(\cache_tag[5][18] ), .op(n7731) );
  nand2_1 U7781 ( .ip1(n10941), .ip2(\cache_tag[11][18] ), .op(n7730) );
  nand2_1 U7782 ( .ip1(n10939), .ip2(\cache_tag[12][18] ), .op(n7729) );
  nand4_1 U7783 ( .ip1(n7732), .ip2(n7731), .ip3(n7730), .ip4(n7729), .op(
        n7748) );
  nand2_1 U7784 ( .ip1(n10931), .ip2(\cache_tag[3][18] ), .op(n7736) );
  nand2_1 U7785 ( .ip1(n10930), .ip2(\cache_tag[1][18] ), .op(n7735) );
  nand2_1 U7786 ( .ip1(n10924), .ip2(\cache_tag[6][18] ), .op(n7734) );
  nand2_1 U7787 ( .ip1(n10932), .ip2(\cache_tag[8][18] ), .op(n7733) );
  nand4_1 U7788 ( .ip1(n7736), .ip2(n7735), .ip3(n7734), .ip4(n7733), .op(
        n7747) );
  nand2_1 U7789 ( .ip1(n10925), .ip2(\cache_tag[2][18] ), .op(n7740) );
  nand2_1 U7790 ( .ip1(n10946), .ip2(\cache_tag[0][18] ), .op(n7739) );
  nand2_1 U7791 ( .ip1(n10923), .ip2(\cache_tag[9][18] ), .op(n7738) );
  nand2_1 U7792 ( .ip1(n10949), .ip2(\cache_tag[13][18] ), .op(n7737) );
  nand4_1 U7793 ( .ip1(n7740), .ip2(n7739), .ip3(n7738), .ip4(n7737), .op(
        n7746) );
  nand2_1 U7794 ( .ip1(n10948), .ip2(\cache_tag[4][18] ), .op(n7744) );
  nand2_1 U7795 ( .ip1(n10922), .ip2(\cache_tag[10][18] ), .op(n7743) );
  nand2_1 U7796 ( .ip1(n10940), .ip2(\cache_tag[15][18] ), .op(n7742) );
  nand2_1 U7797 ( .ip1(n10938), .ip2(\cache_tag[14][18] ), .op(n7741) );
  nand4_1 U7798 ( .ip1(n7744), .ip2(n7743), .ip3(n7742), .ip4(n7741), .op(
        n7745) );
  nor4_1 U7799 ( .ip1(n7748), .ip2(n7747), .ip3(n7746), .ip4(n7745), .op(n7749) );
  xor2_1 U7800 ( .ip1(addr_req[26]), .ip2(n7749), .op(n7750) );
  nand4_1 U7801 ( .ip1(n7752), .ip2(n7751), .ip3(n11358), .ip4(n7750), .op(
        n8110) );
  nand2_1 U7802 ( .ip1(n10925), .ip2(\cache_tag[2][10] ), .op(n7756) );
  nand2_1 U7803 ( .ip1(n10946), .ip2(\cache_tag[0][10] ), .op(n7755) );
  nand2_1 U7804 ( .ip1(n10938), .ip2(\cache_tag[14][10] ), .op(n7754) );
  nand2_1 U7805 ( .ip1(n10932), .ip2(\cache_tag[8][10] ), .op(n7753) );
  nand4_1 U7806 ( .ip1(n7756), .ip2(n7755), .ip3(n7754), .ip4(n7753), .op(
        n7772) );
  nand2_1 U7807 ( .ip1(n10941), .ip2(\cache_tag[11][10] ), .op(n7760) );
  nand2_1 U7808 ( .ip1(n10948), .ip2(\cache_tag[4][10] ), .op(n7759) );
  nand2_1 U7809 ( .ip1(n10931), .ip2(\cache_tag[3][10] ), .op(n7758) );
  nand2_1 U7810 ( .ip1(n10939), .ip2(\cache_tag[12][10] ), .op(n7757) );
  nand4_1 U7811 ( .ip1(n7760), .ip2(n7759), .ip3(n7758), .ip4(n7757), .op(
        n7771) );
  nand2_1 U7812 ( .ip1(n10922), .ip2(\cache_tag[10][10] ), .op(n7764) );
  nand2_1 U7813 ( .ip1(n10923), .ip2(\cache_tag[9][10] ), .op(n7763) );
  nand2_1 U7814 ( .ip1(n10924), .ip2(\cache_tag[6][10] ), .op(n7762) );
  nand2_1 U7815 ( .ip1(n10949), .ip2(\cache_tag[13][10] ), .op(n7761) );
  nand4_1 U7816 ( .ip1(n7764), .ip2(n7763), .ip3(n7762), .ip4(n7761), .op(
        n7770) );
  nand2_1 U7817 ( .ip1(n10933), .ip2(\cache_tag[7][10] ), .op(n7768) );
  nand2_1 U7818 ( .ip1(n10940), .ip2(\cache_tag[15][10] ), .op(n7767) );
  nand2_1 U7819 ( .ip1(n10947), .ip2(\cache_tag[5][10] ), .op(n7766) );
  nand2_1 U7820 ( .ip1(n10930), .ip2(\cache_tag[1][10] ), .op(n7765) );
  nand4_1 U7821 ( .ip1(n7768), .ip2(n7767), .ip3(n7766), .ip4(n7765), .op(
        n7769) );
  nor4_1 U7822 ( .ip1(n7772), .ip2(n7771), .ip3(n7770), .ip4(n7769), .op(n7773) );
  xor2_1 U7823 ( .ip1(addr_req[18]), .ip2(n7773), .op(n7840) );
  nand2_1 U7824 ( .ip1(n10922), .ip2(\cache_tag[10][2] ), .op(n7777) );
  nand2_1 U7825 ( .ip1(n10931), .ip2(\cache_tag[3][2] ), .op(n7776) );
  nand2_1 U7826 ( .ip1(n10925), .ip2(\cache_tag[2][2] ), .op(n7775) );
  nand2_1 U7827 ( .ip1(n10948), .ip2(\cache_tag[4][2] ), .op(n7774) );
  nand4_1 U7828 ( .ip1(n7777), .ip2(n7776), .ip3(n7775), .ip4(n7774), .op(
        n7793) );
  nand2_1 U7829 ( .ip1(n10949), .ip2(\cache_tag[13][2] ), .op(n7781) );
  nand2_1 U7830 ( .ip1(n10933), .ip2(\cache_tag[7][2] ), .op(n7780) );
  nand2_1 U7831 ( .ip1(n10932), .ip2(\cache_tag[8][2] ), .op(n7779) );
  nand2_1 U7832 ( .ip1(n10947), .ip2(\cache_tag[5][2] ), .op(n7778) );
  nand4_1 U7833 ( .ip1(n7781), .ip2(n7780), .ip3(n7779), .ip4(n7778), .op(
        n7792) );
  nand2_1 U7834 ( .ip1(n10930), .ip2(\cache_tag[1][2] ), .op(n7785) );
  nand2_1 U7835 ( .ip1(n10923), .ip2(\cache_tag[9][2] ), .op(n7784) );
  nand2_1 U7836 ( .ip1(n10940), .ip2(\cache_tag[15][2] ), .op(n7783) );
  nand2_1 U7837 ( .ip1(n10946), .ip2(\cache_tag[0][2] ), .op(n7782) );
  nand4_1 U7838 ( .ip1(n7785), .ip2(n7784), .ip3(n7783), .ip4(n7782), .op(
        n7791) );
  nand2_1 U7839 ( .ip1(n10924), .ip2(\cache_tag[6][2] ), .op(n7789) );
  nand2_1 U7840 ( .ip1(n10941), .ip2(\cache_tag[11][2] ), .op(n7788) );
  nand2_1 U7841 ( .ip1(n10938), .ip2(\cache_tag[14][2] ), .op(n7787) );
  nand2_1 U7842 ( .ip1(n10939), .ip2(\cache_tag[12][2] ), .op(n7786) );
  nand4_1 U7843 ( .ip1(n7789), .ip2(n7788), .ip3(n7787), .ip4(n7786), .op(
        n7790) );
  nor4_1 U7844 ( .ip1(n7793), .ip2(n7792), .ip3(n7791), .ip4(n7790), .op(n7794) );
  xor2_1 U7845 ( .ip1(addr_req[10]), .ip2(n7794), .op(n7839) );
  nand2_1 U7846 ( .ip1(n10922), .ip2(\cache_tag[10][23] ), .op(n7798) );
  nand2_1 U7847 ( .ip1(n10925), .ip2(\cache_tag[2][23] ), .op(n7797) );
  nand2_1 U7848 ( .ip1(n10923), .ip2(\cache_tag[9][23] ), .op(n7796) );
  nand2_1 U7849 ( .ip1(n10938), .ip2(\cache_tag[14][23] ), .op(n7795) );
  nand4_1 U7850 ( .ip1(n7798), .ip2(n7797), .ip3(n7796), .ip4(n7795), .op(
        n7814) );
  nand2_1 U7851 ( .ip1(n10947), .ip2(\cache_tag[5][23] ), .op(n7802) );
  nand2_1 U7852 ( .ip1(n10933), .ip2(\cache_tag[7][23] ), .op(n7801) );
  nand2_1 U7853 ( .ip1(n10949), .ip2(\cache_tag[13][23] ), .op(n7800) );
  nand2_1 U7854 ( .ip1(n10932), .ip2(\cache_tag[8][23] ), .op(n7799) );
  nand4_1 U7855 ( .ip1(n7802), .ip2(n7801), .ip3(n7800), .ip4(n7799), .op(
        n7813) );
  nand2_1 U7856 ( .ip1(n10946), .ip2(\cache_tag[0][23] ), .op(n7806) );
  nand2_1 U7857 ( .ip1(n10940), .ip2(\cache_tag[15][23] ), .op(n7805) );
  nand2_1 U7858 ( .ip1(n10930), .ip2(\cache_tag[1][23] ), .op(n7804) );
  nand2_1 U7859 ( .ip1(n10948), .ip2(\cache_tag[4][23] ), .op(n7803) );
  nand4_1 U7860 ( .ip1(n7806), .ip2(n7805), .ip3(n7804), .ip4(n7803), .op(
        n7812) );
  nand2_1 U7861 ( .ip1(n10931), .ip2(\cache_tag[3][23] ), .op(n7810) );
  nand2_1 U7862 ( .ip1(n10924), .ip2(\cache_tag[6][23] ), .op(n7809) );
  nand2_1 U7863 ( .ip1(n10939), .ip2(\cache_tag[12][23] ), .op(n7808) );
  nand2_1 U7864 ( .ip1(n10941), .ip2(\cache_tag[11][23] ), .op(n7807) );
  nand4_1 U7865 ( .ip1(n7810), .ip2(n7809), .ip3(n7808), .ip4(n7807), .op(
        n7811) );
  nor4_1 U7866 ( .ip1(n7814), .ip2(n7813), .ip3(n7812), .ip4(n7811), .op(n7815) );
  xor2_1 U7867 ( .ip1(addr_req[31]), .ip2(n7815), .op(n7838) );
  nand2_1 U7868 ( .ip1(n10923), .ip2(\cache_tag[9][16] ), .op(n7819) );
  nand2_1 U7869 ( .ip1(n10932), .ip2(\cache_tag[8][16] ), .op(n7818) );
  nand2_1 U7870 ( .ip1(n10924), .ip2(\cache_tag[6][16] ), .op(n7817) );
  nand2_1 U7871 ( .ip1(n10946), .ip2(\cache_tag[0][16] ), .op(n7816) );
  nand4_1 U7872 ( .ip1(n7819), .ip2(n7818), .ip3(n7817), .ip4(n7816), .op(
        n7835) );
  nand2_1 U7873 ( .ip1(n10947), .ip2(\cache_tag[5][16] ), .op(n7823) );
  nand2_1 U7874 ( .ip1(n10940), .ip2(\cache_tag[15][16] ), .op(n7822) );
  nand2_1 U7875 ( .ip1(n10922), .ip2(\cache_tag[10][16] ), .op(n7821) );
  nand2_1 U7876 ( .ip1(n10925), .ip2(\cache_tag[2][16] ), .op(n7820) );
  nand4_1 U7877 ( .ip1(n7823), .ip2(n7822), .ip3(n7821), .ip4(n7820), .op(
        n7834) );
  nand2_1 U7878 ( .ip1(n10939), .ip2(\cache_tag[12][16] ), .op(n7827) );
  nand2_1 U7879 ( .ip1(n10941), .ip2(\cache_tag[11][16] ), .op(n7826) );
  nand2_1 U7880 ( .ip1(n10948), .ip2(\cache_tag[4][16] ), .op(n7825) );
  nand2_1 U7881 ( .ip1(n10933), .ip2(\cache_tag[7][16] ), .op(n7824) );
  nand4_1 U7882 ( .ip1(n7827), .ip2(n7826), .ip3(n7825), .ip4(n7824), .op(
        n7833) );
  nand2_1 U7883 ( .ip1(n10949), .ip2(\cache_tag[13][16] ), .op(n7831) );
  nand2_1 U7884 ( .ip1(n10931), .ip2(\cache_tag[3][16] ), .op(n7830) );
  nand2_1 U7885 ( .ip1(n10930), .ip2(\cache_tag[1][16] ), .op(n7829) );
  nand2_1 U7886 ( .ip1(n10938), .ip2(\cache_tag[14][16] ), .op(n7828) );
  nand4_1 U7887 ( .ip1(n7831), .ip2(n7830), .ip3(n7829), .ip4(n7828), .op(
        n7832) );
  nor4_1 U7888 ( .ip1(n7835), .ip2(n7834), .ip3(n7833), .ip4(n7832), .op(n7836) );
  xor2_1 U7889 ( .ip1(addr_req[24]), .ip2(n7836), .op(n7837) );
  nand4_1 U7890 ( .ip1(n7840), .ip2(n7839), .ip3(n7838), .ip4(n7837), .op(
        n8108) );
  nand2_1 U7891 ( .ip1(n10940), .ip2(\cache_tag[15][8] ), .op(n7844) );
  nand2_1 U7892 ( .ip1(n10949), .ip2(\cache_tag[13][8] ), .op(n7843) );
  nand2_1 U7893 ( .ip1(n10923), .ip2(\cache_tag[9][8] ), .op(n7842) );
  nand2_1 U7894 ( .ip1(n10946), .ip2(\cache_tag[0][8] ), .op(n7841) );
  nand4_1 U7895 ( .ip1(n7844), .ip2(n7843), .ip3(n7842), .ip4(n7841), .op(
        n7860) );
  nand2_1 U7896 ( .ip1(n10931), .ip2(\cache_tag[3][8] ), .op(n7848) );
  nand2_1 U7897 ( .ip1(n10930), .ip2(\cache_tag[1][8] ), .op(n7847) );
  nand2_1 U7898 ( .ip1(n10925), .ip2(\cache_tag[2][8] ), .op(n7846) );
  nand2_1 U7899 ( .ip1(n10938), .ip2(\cache_tag[14][8] ), .op(n7845) );
  nand4_1 U7900 ( .ip1(n7848), .ip2(n7847), .ip3(n7846), .ip4(n7845), .op(
        n7859) );
  nand2_1 U7901 ( .ip1(n10924), .ip2(\cache_tag[6][8] ), .op(n7852) );
  nand2_1 U7902 ( .ip1(n10933), .ip2(\cache_tag[7][8] ), .op(n7851) );
  nand2_1 U7903 ( .ip1(n10932), .ip2(\cache_tag[8][8] ), .op(n7850) );
  nand2_1 U7904 ( .ip1(n10939), .ip2(\cache_tag[12][8] ), .op(n7849) );
  nand4_1 U7905 ( .ip1(n7852), .ip2(n7851), .ip3(n7850), .ip4(n7849), .op(
        n7858) );
  nand2_1 U7906 ( .ip1(n10948), .ip2(\cache_tag[4][8] ), .op(n7856) );
  nand2_1 U7907 ( .ip1(n10941), .ip2(\cache_tag[11][8] ), .op(n7855) );
  nand2_1 U7908 ( .ip1(n10922), .ip2(\cache_tag[10][8] ), .op(n7854) );
  nand2_1 U7909 ( .ip1(n10947), .ip2(\cache_tag[5][8] ), .op(n7853) );
  nand4_1 U7910 ( .ip1(n7856), .ip2(n7855), .ip3(n7854), .ip4(n7853), .op(
        n7857) );
  nor4_1 U7911 ( .ip1(n7860), .ip2(n7859), .ip3(n7858), .ip4(n7857), .op(n7861) );
  xor2_1 U7912 ( .ip1(addr_req[16]), .ip2(n7861), .op(n7928) );
  nand2_1 U7913 ( .ip1(n10938), .ip2(\cache_tag[14][3] ), .op(n7865) );
  nand2_1 U7914 ( .ip1(n10924), .ip2(\cache_tag[6][3] ), .op(n7864) );
  nand2_1 U7915 ( .ip1(n10947), .ip2(\cache_tag[5][3] ), .op(n7863) );
  nand2_1 U7916 ( .ip1(n10925), .ip2(\cache_tag[2][3] ), .op(n7862) );
  nand4_1 U7917 ( .ip1(n7865), .ip2(n7864), .ip3(n7863), .ip4(n7862), .op(
        n7881) );
  nand2_1 U7918 ( .ip1(n10940), .ip2(\cache_tag[15][3] ), .op(n7869) );
  nand2_1 U7919 ( .ip1(n10941), .ip2(\cache_tag[11][3] ), .op(n7868) );
  nand2_1 U7920 ( .ip1(n10923), .ip2(\cache_tag[9][3] ), .op(n7867) );
  nand2_1 U7921 ( .ip1(n10949), .ip2(\cache_tag[13][3] ), .op(n7866) );
  nand4_1 U7922 ( .ip1(n7869), .ip2(n7868), .ip3(n7867), .ip4(n7866), .op(
        n7880) );
  nand2_1 U7923 ( .ip1(n10931), .ip2(\cache_tag[3][3] ), .op(n7873) );
  nand2_1 U7924 ( .ip1(n10932), .ip2(\cache_tag[8][3] ), .op(n7872) );
  nand2_1 U7925 ( .ip1(n10933), .ip2(\cache_tag[7][3] ), .op(n7871) );
  nand2_1 U7926 ( .ip1(n10948), .ip2(\cache_tag[4][3] ), .op(n7870) );
  nand4_1 U7927 ( .ip1(n7873), .ip2(n7872), .ip3(n7871), .ip4(n7870), .op(
        n7879) );
  nand2_1 U7928 ( .ip1(n10939), .ip2(\cache_tag[12][3] ), .op(n7877) );
  nand2_1 U7929 ( .ip1(n10930), .ip2(\cache_tag[1][3] ), .op(n7876) );
  nand2_1 U7930 ( .ip1(n10946), .ip2(\cache_tag[0][3] ), .op(n7875) );
  nand2_1 U7931 ( .ip1(n10922), .ip2(\cache_tag[10][3] ), .op(n7874) );
  nand4_1 U7932 ( .ip1(n7877), .ip2(n7876), .ip3(n7875), .ip4(n7874), .op(
        n7878) );
  nor4_1 U7933 ( .ip1(n7881), .ip2(n7880), .ip3(n7879), .ip4(n7878), .op(n7882) );
  xor2_1 U7934 ( .ip1(addr_req[11]), .ip2(n7882), .op(n7927) );
  nand2_1 U7935 ( .ip1(n10946), .ip2(\cache_tag[0][6] ), .op(n7886) );
  nand2_1 U7936 ( .ip1(n10940), .ip2(\cache_tag[15][6] ), .op(n7885) );
  nand2_1 U7937 ( .ip1(n10947), .ip2(\cache_tag[5][6] ), .op(n7884) );
  nand2_1 U7938 ( .ip1(n10924), .ip2(\cache_tag[6][6] ), .op(n7883) );
  nand4_1 U7939 ( .ip1(n7886), .ip2(n7885), .ip3(n7884), .ip4(n7883), .op(
        n7902) );
  nand2_1 U7940 ( .ip1(n10932), .ip2(\cache_tag[8][6] ), .op(n7890) );
  nand2_1 U7941 ( .ip1(n10949), .ip2(\cache_tag[13][6] ), .op(n7889) );
  nand2_1 U7942 ( .ip1(n10948), .ip2(\cache_tag[4][6] ), .op(n7888) );
  nand2_1 U7943 ( .ip1(n10922), .ip2(\cache_tag[10][6] ), .op(n7887) );
  nand4_1 U7944 ( .ip1(n7890), .ip2(n7889), .ip3(n7888), .ip4(n7887), .op(
        n7901) );
  nand2_1 U7945 ( .ip1(n10931), .ip2(\cache_tag[3][6] ), .op(n7894) );
  nand2_1 U7946 ( .ip1(n10923), .ip2(\cache_tag[9][6] ), .op(n7893) );
  nand2_1 U7947 ( .ip1(n10939), .ip2(\cache_tag[12][6] ), .op(n7892) );
  nand2_1 U7948 ( .ip1(n10930), .ip2(\cache_tag[1][6] ), .op(n7891) );
  nand4_1 U7949 ( .ip1(n7894), .ip2(n7893), .ip3(n7892), .ip4(n7891), .op(
        n7900) );
  nand2_1 U7950 ( .ip1(n10933), .ip2(\cache_tag[7][6] ), .op(n7898) );
  nand2_1 U7951 ( .ip1(n10941), .ip2(\cache_tag[11][6] ), .op(n7897) );
  nand2_1 U7952 ( .ip1(n10938), .ip2(\cache_tag[14][6] ), .op(n7896) );
  nand2_1 U7953 ( .ip1(n10925), .ip2(\cache_tag[2][6] ), .op(n7895) );
  nand4_1 U7954 ( .ip1(n7898), .ip2(n7897), .ip3(n7896), .ip4(n7895), .op(
        n7899) );
  nor4_1 U7955 ( .ip1(n7902), .ip2(n7901), .ip3(n7900), .ip4(n7899), .op(n7903) );
  xor2_1 U7956 ( .ip1(addr_req[14]), .ip2(n7903), .op(n7926) );
  nand2_1 U7957 ( .ip1(n10940), .ip2(\cache_tag[15][19] ), .op(n7907) );
  nand2_1 U7958 ( .ip1(n10938), .ip2(\cache_tag[14][19] ), .op(n7906) );
  nand2_1 U7959 ( .ip1(n10947), .ip2(\cache_tag[5][19] ), .op(n7905) );
  nand2_1 U7960 ( .ip1(n10941), .ip2(\cache_tag[11][19] ), .op(n7904) );
  nand4_1 U7961 ( .ip1(n7907), .ip2(n7906), .ip3(n7905), .ip4(n7904), .op(
        n7923) );
  nand2_1 U7962 ( .ip1(n10923), .ip2(\cache_tag[9][19] ), .op(n7911) );
  nand2_1 U7963 ( .ip1(n10949), .ip2(\cache_tag[13][19] ), .op(n7910) );
  nand2_1 U7964 ( .ip1(n10930), .ip2(\cache_tag[1][19] ), .op(n7909) );
  nand2_1 U7965 ( .ip1(n10932), .ip2(\cache_tag[8][19] ), .op(n7908) );
  nand4_1 U7966 ( .ip1(n7911), .ip2(n7910), .ip3(n7909), .ip4(n7908), .op(
        n7922) );
  nand2_1 U7967 ( .ip1(n10939), .ip2(\cache_tag[12][19] ), .op(n7915) );
  nand2_1 U7968 ( .ip1(n10948), .ip2(\cache_tag[4][19] ), .op(n7914) );
  nand2_1 U7969 ( .ip1(n10924), .ip2(\cache_tag[6][19] ), .op(n7913) );
  nand2_1 U7970 ( .ip1(n10946), .ip2(\cache_tag[0][19] ), .op(n7912) );
  nand4_1 U7971 ( .ip1(n7915), .ip2(n7914), .ip3(n7913), .ip4(n7912), .op(
        n7921) );
  nand2_1 U7972 ( .ip1(n10925), .ip2(\cache_tag[2][19] ), .op(n7919) );
  nand2_1 U7973 ( .ip1(n10931), .ip2(\cache_tag[3][19] ), .op(n7918) );
  nand2_1 U7974 ( .ip1(n10922), .ip2(\cache_tag[10][19] ), .op(n7917) );
  nand2_1 U7975 ( .ip1(n10933), .ip2(\cache_tag[7][19] ), .op(n7916) );
  nand4_1 U7976 ( .ip1(n7919), .ip2(n7918), .ip3(n7917), .ip4(n7916), .op(
        n7920) );
  nor4_1 U7977 ( .ip1(n7923), .ip2(n7922), .ip3(n7921), .ip4(n7920), .op(n7924) );
  xor2_1 U7978 ( .ip1(addr_req[27]), .ip2(n7924), .op(n7925) );
  nand4_1 U7979 ( .ip1(n7928), .ip2(n7927), .ip3(n7926), .ip4(n7925), .op(
        n8107) );
  nand2_1 U7980 ( .ip1(n10931), .ip2(\cache_tag[3][21] ), .op(n7932) );
  nand2_1 U7981 ( .ip1(n10924), .ip2(\cache_tag[6][21] ), .op(n7931) );
  nand2_1 U7982 ( .ip1(n10948), .ip2(\cache_tag[4][21] ), .op(n7930) );
  nand2_1 U7983 ( .ip1(n10941), .ip2(\cache_tag[11][21] ), .op(n7929) );
  nand4_1 U7984 ( .ip1(n7932), .ip2(n7931), .ip3(n7930), .ip4(n7929), .op(
        n7948) );
  nand2_1 U7985 ( .ip1(n10938), .ip2(\cache_tag[14][21] ), .op(n7936) );
  nand2_1 U7986 ( .ip1(n10930), .ip2(\cache_tag[1][21] ), .op(n7935) );
  nand2_1 U7987 ( .ip1(n10949), .ip2(\cache_tag[13][21] ), .op(n7934) );
  nand2_1 U7988 ( .ip1(n10925), .ip2(\cache_tag[2][21] ), .op(n7933) );
  nand4_1 U7989 ( .ip1(n7936), .ip2(n7935), .ip3(n7934), .ip4(n7933), .op(
        n7947) );
  nand2_1 U7990 ( .ip1(n10932), .ip2(\cache_tag[8][21] ), .op(n7940) );
  nand2_1 U7991 ( .ip1(n10940), .ip2(\cache_tag[15][21] ), .op(n7939) );
  nand2_1 U7992 ( .ip1(n10933), .ip2(\cache_tag[7][21] ), .op(n7938) );
  nand2_1 U7993 ( .ip1(n10923), .ip2(\cache_tag[9][21] ), .op(n7937) );
  nand4_1 U7994 ( .ip1(n7940), .ip2(n7939), .ip3(n7938), .ip4(n7937), .op(
        n7946) );
  nand2_1 U7995 ( .ip1(n10922), .ip2(\cache_tag[10][21] ), .op(n7944) );
  nand2_1 U7996 ( .ip1(n10947), .ip2(\cache_tag[5][21] ), .op(n7943) );
  nand2_1 U7997 ( .ip1(n10939), .ip2(\cache_tag[12][21] ), .op(n7942) );
  nand2_1 U7998 ( .ip1(n10946), .ip2(\cache_tag[0][21] ), .op(n7941) );
  nand4_1 U7999 ( .ip1(n7944), .ip2(n7943), .ip3(n7942), .ip4(n7941), .op(
        n7945) );
  nor4_1 U8000 ( .ip1(n7948), .ip2(n7947), .ip3(n7946), .ip4(n7945), .op(n7949) );
  xor2_1 U8001 ( .ip1(addr_req[29]), .ip2(n7949), .op(n8016) );
  nand2_1 U8002 ( .ip1(n10930), .ip2(\cache_tag[1][0] ), .op(n7953) );
  nand2_1 U8003 ( .ip1(n10940), .ip2(\cache_tag[15][0] ), .op(n7952) );
  nand2_1 U8004 ( .ip1(n10924), .ip2(\cache_tag[6][0] ), .op(n7951) );
  nand2_1 U8005 ( .ip1(n10941), .ip2(\cache_tag[11][0] ), .op(n7950) );
  nand4_1 U8006 ( .ip1(n7953), .ip2(n7952), .ip3(n7951), .ip4(n7950), .op(
        n7969) );
  nand2_1 U8007 ( .ip1(n10923), .ip2(\cache_tag[9][0] ), .op(n7957) );
  nand2_1 U8008 ( .ip1(n10938), .ip2(\cache_tag[14][0] ), .op(n7956) );
  nand2_1 U8009 ( .ip1(n10931), .ip2(\cache_tag[3][0] ), .op(n7955) );
  nand2_1 U8010 ( .ip1(n10939), .ip2(\cache_tag[12][0] ), .op(n7954) );
  nand4_1 U8011 ( .ip1(n7957), .ip2(n7956), .ip3(n7955), .ip4(n7954), .op(
        n7968) );
  nand2_1 U8012 ( .ip1(n10922), .ip2(\cache_tag[10][0] ), .op(n7961) );
  nand2_1 U8013 ( .ip1(n10949), .ip2(\cache_tag[13][0] ), .op(n7960) );
  nand2_1 U8014 ( .ip1(n10948), .ip2(\cache_tag[4][0] ), .op(n7959) );
  nand2_1 U8015 ( .ip1(n10947), .ip2(\cache_tag[5][0] ), .op(n7958) );
  nand4_1 U8016 ( .ip1(n7961), .ip2(n7960), .ip3(n7959), .ip4(n7958), .op(
        n7967) );
  nand2_1 U8017 ( .ip1(n10925), .ip2(\cache_tag[2][0] ), .op(n7965) );
  nand2_1 U8018 ( .ip1(n10932), .ip2(\cache_tag[8][0] ), .op(n7964) );
  nand2_1 U8019 ( .ip1(n10946), .ip2(\cache_tag[0][0] ), .op(n7963) );
  nand2_1 U8020 ( .ip1(n10933), .ip2(\cache_tag[7][0] ), .op(n7962) );
  nand4_1 U8021 ( .ip1(n7965), .ip2(n7964), .ip3(n7963), .ip4(n7962), .op(
        n7966) );
  nor4_1 U8022 ( .ip1(n7969), .ip2(n7968), .ip3(n7967), .ip4(n7966), .op(n7970) );
  xor2_1 U8023 ( .ip1(addr_req[8]), .ip2(n7970), .op(n8015) );
  nand2_1 U8024 ( .ip1(n10931), .ip2(\cache_tag[3][7] ), .op(n7974) );
  nand2_1 U8025 ( .ip1(n10939), .ip2(\cache_tag[12][7] ), .op(n7973) );
  nand2_1 U8026 ( .ip1(n10948), .ip2(\cache_tag[4][7] ), .op(n7972) );
  nand2_1 U8027 ( .ip1(n10933), .ip2(\cache_tag[7][7] ), .op(n7971) );
  nand4_1 U8028 ( .ip1(n7974), .ip2(n7973), .ip3(n7972), .ip4(n7971), .op(
        n7990) );
  nand2_1 U8029 ( .ip1(n10946), .ip2(\cache_tag[0][7] ), .op(n7978) );
  nand2_1 U8030 ( .ip1(n10922), .ip2(\cache_tag[10][7] ), .op(n7977) );
  nand2_1 U8031 ( .ip1(n10924), .ip2(\cache_tag[6][7] ), .op(n7976) );
  nand2_1 U8032 ( .ip1(n10941), .ip2(\cache_tag[11][7] ), .op(n7975) );
  nand4_1 U8033 ( .ip1(n7978), .ip2(n7977), .ip3(n7976), .ip4(n7975), .op(
        n7989) );
  nand2_1 U8034 ( .ip1(n10932), .ip2(\cache_tag[8][7] ), .op(n7982) );
  nand2_1 U8035 ( .ip1(n10923), .ip2(\cache_tag[9][7] ), .op(n7981) );
  nand2_1 U8036 ( .ip1(n10930), .ip2(\cache_tag[1][7] ), .op(n7980) );
  nand2_1 U8037 ( .ip1(n10949), .ip2(\cache_tag[13][7] ), .op(n7979) );
  nand4_1 U8038 ( .ip1(n7982), .ip2(n7981), .ip3(n7980), .ip4(n7979), .op(
        n7988) );
  nand2_1 U8039 ( .ip1(n10925), .ip2(\cache_tag[2][7] ), .op(n7986) );
  nand2_1 U8040 ( .ip1(n10947), .ip2(\cache_tag[5][7] ), .op(n7985) );
  nand2_1 U8041 ( .ip1(n10938), .ip2(\cache_tag[14][7] ), .op(n7984) );
  nand2_1 U8042 ( .ip1(n10940), .ip2(\cache_tag[15][7] ), .op(n7983) );
  nand4_1 U8043 ( .ip1(n7986), .ip2(n7985), .ip3(n7984), .ip4(n7983), .op(
        n7987) );
  nor4_1 U8044 ( .ip1(n7990), .ip2(n7989), .ip3(n7988), .ip4(n7987), .op(n7991) );
  xor2_1 U8045 ( .ip1(addr_req[15]), .ip2(n7991), .op(n8014) );
  nand2_1 U8046 ( .ip1(n10925), .ip2(\cache_tag[2][22] ), .op(n7995) );
  nand2_1 U8047 ( .ip1(n10940), .ip2(\cache_tag[15][22] ), .op(n7994) );
  nand2_1 U8048 ( .ip1(n10949), .ip2(\cache_tag[13][22] ), .op(n7993) );
  nand2_1 U8049 ( .ip1(n10932), .ip2(\cache_tag[8][22] ), .op(n7992) );
  nand4_1 U8050 ( .ip1(n7995), .ip2(n7994), .ip3(n7993), .ip4(n7992), .op(
        n8011) );
  nand2_1 U8051 ( .ip1(n10931), .ip2(\cache_tag[3][22] ), .op(n7999) );
  nand2_1 U8052 ( .ip1(n10930), .ip2(\cache_tag[1][22] ), .op(n7998) );
  nand2_1 U8053 ( .ip1(n10922), .ip2(\cache_tag[10][22] ), .op(n7997) );
  nand2_1 U8054 ( .ip1(n10933), .ip2(\cache_tag[7][22] ), .op(n7996) );
  nand4_1 U8055 ( .ip1(n7999), .ip2(n7998), .ip3(n7997), .ip4(n7996), .op(
        n8010) );
  nand2_1 U8056 ( .ip1(n10923), .ip2(\cache_tag[9][22] ), .op(n8003) );
  nand2_1 U8057 ( .ip1(n10924), .ip2(\cache_tag[6][22] ), .op(n8002) );
  nand2_1 U8058 ( .ip1(n10946), .ip2(\cache_tag[0][22] ), .op(n8001) );
  nand2_1 U8059 ( .ip1(n10947), .ip2(\cache_tag[5][22] ), .op(n8000) );
  nand4_1 U8060 ( .ip1(n8003), .ip2(n8002), .ip3(n8001), .ip4(n8000), .op(
        n8009) );
  nand2_1 U8061 ( .ip1(n10938), .ip2(\cache_tag[14][22] ), .op(n8007) );
  nand2_1 U8062 ( .ip1(n10939), .ip2(\cache_tag[12][22] ), .op(n8006) );
  nand2_1 U8063 ( .ip1(n10941), .ip2(\cache_tag[11][22] ), .op(n8005) );
  nand2_1 U8064 ( .ip1(n10948), .ip2(\cache_tag[4][22] ), .op(n8004) );
  nand4_1 U8065 ( .ip1(n8007), .ip2(n8006), .ip3(n8005), .ip4(n8004), .op(
        n8008) );
  nor4_1 U8066 ( .ip1(n8011), .ip2(n8010), .ip3(n8009), .ip4(n8008), .op(n8012) );
  xor2_1 U8067 ( .ip1(addr_req[30]), .ip2(n8012), .op(n8013) );
  nand4_1 U8068 ( .ip1(n8016), .ip2(n8015), .ip3(n8014), .ip4(n8013), .op(
        n8106) );
  nand2_1 U8069 ( .ip1(n10922), .ip2(\cache_tag[10][5] ), .op(n8020) );
  nand2_1 U8070 ( .ip1(n10938), .ip2(\cache_tag[14][5] ), .op(n8019) );
  nand2_1 U8071 ( .ip1(n10941), .ip2(\cache_tag[11][5] ), .op(n8018) );
  nand2_1 U8072 ( .ip1(n10923), .ip2(\cache_tag[9][5] ), .op(n8017) );
  nand4_1 U8073 ( .ip1(n8020), .ip2(n8019), .ip3(n8018), .ip4(n8017), .op(
        n8036) );
  nand2_1 U8074 ( .ip1(n10930), .ip2(\cache_tag[1][5] ), .op(n8024) );
  nand2_1 U8075 ( .ip1(n10940), .ip2(\cache_tag[15][5] ), .op(n8023) );
  nand2_1 U8076 ( .ip1(n10932), .ip2(\cache_tag[8][5] ), .op(n8022) );
  nand2_1 U8077 ( .ip1(n10925), .ip2(\cache_tag[2][5] ), .op(n8021) );
  nand4_1 U8078 ( .ip1(n8024), .ip2(n8023), .ip3(n8022), .ip4(n8021), .op(
        n8035) );
  nand2_1 U8079 ( .ip1(n10947), .ip2(\cache_tag[5][5] ), .op(n8028) );
  nand2_1 U8080 ( .ip1(n10948), .ip2(\cache_tag[4][5] ), .op(n8027) );
  nand2_1 U8081 ( .ip1(n10931), .ip2(\cache_tag[3][5] ), .op(n8026) );
  nand2_1 U8082 ( .ip1(n10933), .ip2(\cache_tag[7][5] ), .op(n8025) );
  nand4_1 U8083 ( .ip1(n8028), .ip2(n8027), .ip3(n8026), .ip4(n8025), .op(
        n8034) );
  nand2_1 U8084 ( .ip1(n10949), .ip2(\cache_tag[13][5] ), .op(n8032) );
  nand2_1 U8085 ( .ip1(n10939), .ip2(\cache_tag[12][5] ), .op(n8031) );
  nand2_1 U8086 ( .ip1(n10924), .ip2(\cache_tag[6][5] ), .op(n8030) );
  nand2_1 U8087 ( .ip1(n10946), .ip2(\cache_tag[0][5] ), .op(n8029) );
  nand4_1 U8088 ( .ip1(n8032), .ip2(n8031), .ip3(n8030), .ip4(n8029), .op(
        n8033) );
  nor4_1 U8089 ( .ip1(n8036), .ip2(n8035), .ip3(n8034), .ip4(n8033), .op(n8037) );
  xor2_1 U8090 ( .ip1(addr_req[13]), .ip2(n8037), .op(n8104) );
  nand2_1 U8091 ( .ip1(n10941), .ip2(\cache_tag[11][1] ), .op(n8041) );
  nand2_1 U8092 ( .ip1(n10922), .ip2(\cache_tag[10][1] ), .op(n8040) );
  nand2_1 U8093 ( .ip1(n10925), .ip2(\cache_tag[2][1] ), .op(n8039) );
  nand2_1 U8094 ( .ip1(n10946), .ip2(\cache_tag[0][1] ), .op(n8038) );
  nand4_1 U8095 ( .ip1(n8041), .ip2(n8040), .ip3(n8039), .ip4(n8038), .op(
        n8057) );
  nand2_1 U8096 ( .ip1(n10923), .ip2(\cache_tag[9][1] ), .op(n8045) );
  nand2_1 U8097 ( .ip1(n10938), .ip2(\cache_tag[14][1] ), .op(n8044) );
  nand2_1 U8098 ( .ip1(n10948), .ip2(\cache_tag[4][1] ), .op(n8043) );
  nand2_1 U8099 ( .ip1(n10924), .ip2(\cache_tag[6][1] ), .op(n8042) );
  nand4_1 U8100 ( .ip1(n8045), .ip2(n8044), .ip3(n8043), .ip4(n8042), .op(
        n8056) );
  nand2_1 U8101 ( .ip1(n10930), .ip2(\cache_tag[1][1] ), .op(n8049) );
  nand2_1 U8102 ( .ip1(n10940), .ip2(\cache_tag[15][1] ), .op(n8048) );
  nand2_1 U8103 ( .ip1(n10932), .ip2(\cache_tag[8][1] ), .op(n8047) );
  nand2_1 U8104 ( .ip1(n10933), .ip2(\cache_tag[7][1] ), .op(n8046) );
  nand4_1 U8105 ( .ip1(n8049), .ip2(n8048), .ip3(n8047), .ip4(n8046), .op(
        n8055) );
  nand2_1 U8106 ( .ip1(n10947), .ip2(\cache_tag[5][1] ), .op(n8053) );
  nand2_1 U8107 ( .ip1(n10931), .ip2(\cache_tag[3][1] ), .op(n8052) );
  nand2_1 U8108 ( .ip1(n10949), .ip2(\cache_tag[13][1] ), .op(n8051) );
  nand2_1 U8109 ( .ip1(n10939), .ip2(\cache_tag[12][1] ), .op(n8050) );
  nand4_1 U8110 ( .ip1(n8053), .ip2(n8052), .ip3(n8051), .ip4(n8050), .op(
        n8054) );
  nor4_1 U8111 ( .ip1(n8057), .ip2(n8056), .ip3(n8055), .ip4(n8054), .op(n8058) );
  xor2_1 U8112 ( .ip1(addr_req[9]), .ip2(n8058), .op(n8103) );
  nand2_1 U8113 ( .ip1(n10938), .ip2(\cache_tag[14][17] ), .op(n8062) );
  nand2_1 U8114 ( .ip1(n10940), .ip2(\cache_tag[15][17] ), .op(n8061) );
  nand2_1 U8115 ( .ip1(n10941), .ip2(\cache_tag[11][17] ), .op(n8060) );
  nand2_1 U8116 ( .ip1(n10933), .ip2(\cache_tag[7][17] ), .op(n8059) );
  nand4_1 U8117 ( .ip1(n8062), .ip2(n8061), .ip3(n8060), .ip4(n8059), .op(
        n8078) );
  nand2_1 U8118 ( .ip1(n10948), .ip2(\cache_tag[4][17] ), .op(n8066) );
  nand2_1 U8119 ( .ip1(n10946), .ip2(\cache_tag[0][17] ), .op(n8065) );
  nand2_1 U8120 ( .ip1(n10922), .ip2(\cache_tag[10][17] ), .op(n8064) );
  nand2_1 U8121 ( .ip1(n10930), .ip2(\cache_tag[1][17] ), .op(n8063) );
  nand4_1 U8122 ( .ip1(n8066), .ip2(n8065), .ip3(n8064), .ip4(n8063), .op(
        n8077) );
  nand2_1 U8123 ( .ip1(n10923), .ip2(\cache_tag[9][17] ), .op(n8070) );
  nand2_1 U8124 ( .ip1(n10949), .ip2(\cache_tag[13][17] ), .op(n8069) );
  nand2_1 U8125 ( .ip1(n10932), .ip2(\cache_tag[8][17] ), .op(n8068) );
  nand2_1 U8126 ( .ip1(n10924), .ip2(\cache_tag[6][17] ), .op(n8067) );
  nand4_1 U8127 ( .ip1(n8070), .ip2(n8069), .ip3(n8068), .ip4(n8067), .op(
        n8076) );
  nand2_1 U8128 ( .ip1(n10925), .ip2(\cache_tag[2][17] ), .op(n8074) );
  nand2_1 U8129 ( .ip1(n10931), .ip2(\cache_tag[3][17] ), .op(n8073) );
  nand2_1 U8130 ( .ip1(n10939), .ip2(\cache_tag[12][17] ), .op(n8072) );
  nand2_1 U8131 ( .ip1(n10947), .ip2(\cache_tag[5][17] ), .op(n8071) );
  nand4_1 U8132 ( .ip1(n8074), .ip2(n8073), .ip3(n8072), .ip4(n8071), .op(
        n8075) );
  nor4_1 U8133 ( .ip1(n8078), .ip2(n8077), .ip3(n8076), .ip4(n8075), .op(n8079) );
  xor2_1 U8134 ( .ip1(addr_req[25]), .ip2(n8079), .op(n8102) );
  nand2_1 U8135 ( .ip1(n10938), .ip2(\cache_tag[14][4] ), .op(n8083) );
  nand2_1 U8136 ( .ip1(n10948), .ip2(\cache_tag[4][4] ), .op(n8082) );
  nand2_1 U8137 ( .ip1(n10925), .ip2(\cache_tag[2][4] ), .op(n8081) );
  nand2_1 U8138 ( .ip1(n10949), .ip2(\cache_tag[13][4] ), .op(n8080) );
  nand4_1 U8139 ( .ip1(n8083), .ip2(n8082), .ip3(n8081), .ip4(n8080), .op(
        n8099) );
  nand2_1 U8140 ( .ip1(n10931), .ip2(\cache_tag[3][4] ), .op(n8087) );
  nand2_1 U8141 ( .ip1(n10946), .ip2(\cache_tag[0][4] ), .op(n8086) );
  nand2_1 U8142 ( .ip1(n10941), .ip2(\cache_tag[11][4] ), .op(n8085) );
  nand2_1 U8143 ( .ip1(n10940), .ip2(\cache_tag[15][4] ), .op(n8084) );
  nand4_1 U8144 ( .ip1(n8087), .ip2(n8086), .ip3(n8085), .ip4(n8084), .op(
        n8098) );
  nand2_1 U8145 ( .ip1(n10933), .ip2(\cache_tag[7][4] ), .op(n8091) );
  nand2_1 U8146 ( .ip1(n10932), .ip2(\cache_tag[8][4] ), .op(n8090) );
  nand2_1 U8147 ( .ip1(n10924), .ip2(\cache_tag[6][4] ), .op(n8089) );
  nand2_1 U8148 ( .ip1(n10930), .ip2(\cache_tag[1][4] ), .op(n8088) );
  nand4_1 U8149 ( .ip1(n8091), .ip2(n8090), .ip3(n8089), .ip4(n8088), .op(
        n8097) );
  nand2_1 U8150 ( .ip1(n10923), .ip2(\cache_tag[9][4] ), .op(n8095) );
  nand2_1 U8151 ( .ip1(n10947), .ip2(\cache_tag[5][4] ), .op(n8094) );
  nand2_1 U8152 ( .ip1(n10939), .ip2(\cache_tag[12][4] ), .op(n8093) );
  nand2_1 U8153 ( .ip1(n10922), .ip2(\cache_tag[10][4] ), .op(n8092) );
  nand4_1 U8154 ( .ip1(n8095), .ip2(n8094), .ip3(n8093), .ip4(n8092), .op(
        n8096) );
  nor4_1 U8155 ( .ip1(n8099), .ip2(n8098), .ip3(n8097), .ip4(n8096), .op(n8100) );
  xor2_1 U8156 ( .ip1(addr_req[12]), .ip2(n8100), .op(n8101) );
  nand4_1 U8157 ( .ip1(n8104), .ip2(n8103), .ip3(n8102), .ip4(n8101), .op(
        n8105) );
  or4_1 U8158 ( .ip1(n8108), .ip2(n8107), .ip3(n8106), .ip4(n8105), .op(n8109)
         );
  nor4_1 U8159 ( .ip1(n8112), .ip2(n8111), .ip3(n8110), .ip4(n8109), .op(
        n11360) );
  or2_1 U8160 ( .ip1(n8119), .ip2(n11360), .op(n8114) );
  or2_1 U8161 ( .ip1(n11361), .ip2(n11360), .op(n8113) );
  nand2_1 U8162 ( .ip1(n8114), .ip2(n8113), .op(n7412) );
  inv_1 U8163 ( .ip(n8115), .op(n8117) );
  nor4_1 U8164 ( .ip1(state[3]), .ip2(state[1]), .ip3(n8116), .ip4(n8117), 
        .op(n8122) );
  nor4_1 U8165 ( .ip1(state[2]), .ip2(state[1]), .ip3(n8118), .ip4(n8117), 
        .op(n8126) );
  nor2_1 U8166 ( .ip1(n8122), .ip2(n8126), .op(n8132) );
  nor2_1 U8167 ( .ip1(mem_done), .ip2(n8132), .op(n8133) );
  nand2_1 U8168 ( .ip1(state[3]), .ip2(n8133), .op(n8125) );
  or3_1 U8169 ( .ip1(hit), .ip2(n8119), .ip3(dirty), .op(n8120) );
  nand2_1 U8170 ( .ip1(valid), .ip2(n8120), .op(n8121) );
  nand2_1 U8171 ( .ip1(n12287), .ip2(n8121), .op(n8124) );
  nand2_1 U8172 ( .ip1(mem_done), .ip2(n8122), .op(n8123) );
  nand3_1 U8173 ( .ip1(n8125), .ip2(n8124), .ip3(n8123), .op(n12325) );
  nand2_1 U8174 ( .ip1(mem_done), .ip2(n8126), .op(n8129) );
  nand2_1 U8175 ( .ip1(miss), .ip2(dirty), .op(n8127) );
  nand4_1 U8176 ( .ip1(hit), .ip2(n12287), .ip3(valid), .ip4(n8127), .op(n8128) );
  nand2_1 U8177 ( .ip1(n8129), .ip2(n8128), .op(n12323) );
  inv_1 U8178 ( .ip(n12324), .op(n12327) );
  inv_1 U8179 ( .ip(n12324), .op(n12328) );
  inv_1 U8180 ( .ip(n12324), .op(n12329) );
  inv_1 U8181 ( .ip(n12324), .op(n12330) );
  inv_1 U8182 ( .ip(n12324), .op(n12331) );
  inv_1 U8183 ( .ip(n12324), .op(n12332) );
  inv_1 U8184 ( .ip(n12324), .op(n12333) );
  nand3_1 U8186 ( .ip1(n8132), .ip2(n8131), .ip3(n8130), .op(N3691) );
  inv_1 U8187 ( .ip(N3691), .op(next_state[0]) );
  nand2_1 U8188 ( .ip1(state[2]), .ip2(n8133), .op(n8135) );
  nand4_1 U8189 ( .ip1(n12287), .ip2(miss), .ip3(valid), .ip4(dirty), .op(
        n8134) );
  nand2_1 U8190 ( .ip1(n8135), .ip2(n8134), .op(next_state[2]) );
  inv_1 U8191 ( .ip(busy_mem), .op(n10898) );
  nand2_1 U8192 ( .ip1(next_state[2]), .ip2(n10898), .op(n12252) );
  nor2_1 U8193 ( .ip1(n12252), .ip2(n12324), .op(n8211) );
  inv_1 U8194 ( .ip(n8211), .op(n10873) );
  nor3_1 U8195 ( .ip1(mem_data_cnt[3]), .ip2(mem_data_cnt[2]), .ip3(n10873), 
        .op(n10828) );
  inv_1 U8196 ( .ip(addr_resp[5]), .op(n8139) );
  nand2_1 U8197 ( .ip1(addr_resp[6]), .ip2(n8139), .op(n8160) );
  nor3_1 U8198 ( .ip1(addr_resp[7]), .ip2(addr_resp[4]), .ip3(n8160), .op(
        n12201) );
  buf_1 U8199 ( .ip(n12201), .op(n12164) );
  inv_1 U8200 ( .ip(n12164), .op(n8136) );
  inv_1 U8201 ( .ip(n8136), .op(n12243) );
  inv_1 U8202 ( .ip(n8136), .op(n8906) );
  nand2_1 U8203 ( .ip1(n8906), .ip2(\cache_data[4][0] ), .op(n8143) );
  inv_1 U8204 ( .ip(addr_resp[4]), .op(n8138) );
  nand2_1 U8205 ( .ip1(addr_resp[7]), .ip2(n8138), .op(n8162) );
  nor3_1 U8206 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .ip3(n8162), .op(
        n12121) );
  buf_1 U8207 ( .ip(n12121), .op(n12234) );
  inv_1 U8208 ( .ip(n12234), .op(n8137) );
  inv_1 U8209 ( .ip(n8137), .op(n12191) );
  nand2_1 U8210 ( .ip1(n12121), .ip2(\cache_data[8][0] ), .op(n8142) );
  or2_1 U8211 ( .ip1(n8138), .ip2(addr_resp[7]), .op(n8159) );
  or2_1 U8212 ( .ip1(n8139), .ip2(addr_resp[6]), .op(n8158) );
  nor2_1 U8213 ( .ip1(n8159), .ip2(n8158), .op(n12219) );
  inv_1 U8214 ( .ip(n11476), .op(n11317) );
  nand2_1 U8215 ( .ip1(n11317), .ip2(\cache_data[3][0] ), .op(n8141) );
  nor2_1 U8216 ( .ip1(n8160), .ip2(n8162), .op(n12207) );
  buf_1 U8217 ( .ip(n12207), .op(n12030) );
  inv_1 U8218 ( .ip(n11551), .op(n12227) );
  nand2_1 U8219 ( .ip1(n12207), .ip2(\cache_data[12][0] ), .op(n8140) );
  nand4_1 U8220 ( .ip1(n8143), .ip2(n8142), .ip3(n8141), .ip4(n8140), .op(
        n8170) );
  nand2_1 U8221 ( .ip1(addr_resp[7]), .ip2(addr_resp[4]), .op(n8152) );
  nor3_1 U8222 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .ip3(n8152), .op(
        n12126) );
  buf_1 U8223 ( .ip(n12126), .op(n12152) );
  inv_1 U8224 ( .ip(n12152), .op(n8144) );
  inv_1 U8225 ( .ip(n8144), .op(n12241) );
  nand2_1 U8226 ( .ip1(n12126), .ip2(\cache_data[9][0] ), .op(n8150) );
  nor2_1 U8227 ( .ip1(n8160), .ip2(n8152), .op(n12142) );
  buf_1 U8228 ( .ip(n12142), .op(n12242) );
  inv_1 U8229 ( .ip(n12242), .op(n8145) );
  inv_1 U8230 ( .ip(n8145), .op(n12165) );
  inv_1 U8231 ( .ip(n8145), .op(n8899) );
  nand2_1 U8232 ( .ip1(n8899), .ip2(\cache_data[13][0] ), .op(n8149) );
  nor3_1 U8233 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .ip3(n8159), .op(
        n12120) );
  inv_1 U8234 ( .ip(n11459), .op(n8894) );
  nand2_1 U8235 ( .ip1(n8894), .ip2(\cache_data[1][0] ), .op(n8148) );
  nor2_1 U8236 ( .ip1(n8162), .ip2(n8158), .op(n12235) );
  inv_1 U8237 ( .ip(n12235), .op(n8146) );
  inv_1 U8238 ( .ip(n8146), .op(n12196) );
  nand2_1 U8239 ( .ip1(n12196), .ip2(\cache_data[10][0] ), .op(n8147) );
  nand4_1 U8240 ( .ip1(n8150), .ip2(n8149), .ip3(n8148), .ip4(n8147), .op(
        n8169) );
  nand2_1 U8241 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .op(n8161) );
  nor3_1 U8242 ( .ip1(addr_resp[7]), .ip2(addr_resp[4]), .ip3(n8161), .op(
        n12179) );
  buf_1 U8243 ( .ip(n12179), .op(n10305) );
  inv_1 U8244 ( .ip(n11502), .op(n8905) );
  nand2_1 U8245 ( .ip1(n8905), .ip2(\cache_data[6][0] ), .op(n8157) );
  nor2_1 U8246 ( .ip1(n8158), .ip2(n8152), .op(n12096) );
  buf_1 U8247 ( .ip(n12096), .op(n12170) );
  inv_1 U8248 ( .ip(n12170), .op(n8151) );
  inv_1 U8249 ( .ip(n8151), .op(n11927) );
  nand2_1 U8250 ( .ip1(n12096), .ip2(\cache_data[11][0] ), .op(n8156) );
  nor2_1 U8251 ( .ip1(n8152), .ip2(n8161), .op(n12221) );
  buf_1 U8252 ( .ip(n12221), .op(n10975) );
  nand2_1 U8253 ( .ip1(n10975), .ip2(\cache_data[15][0] ), .op(n8155) );
  nor2_1 U8254 ( .ip1(n8159), .ip2(n8161), .op(n12226) );
  buf_1 U8255 ( .ip(n12226), .op(n12143) );
  inv_1 U8256 ( .ip(n12143), .op(n8153) );
  inv_1 U8257 ( .ip(n8153), .op(n12202) );
  nand2_1 U8258 ( .ip1(n12226), .ip2(\cache_data[7][0] ), .op(n8154) );
  nand4_1 U8259 ( .ip1(n8157), .ip2(n8156), .ip3(n8155), .ip4(n8154), .op(
        n8168) );
  nor4_1 U8260 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .ip3(addr_resp[7]), 
        .ip4(addr_resp[4]), .op(n12233) );
  inv_1 U8261 ( .ip(n8923), .op(n8911) );
  nand2_1 U8262 ( .ip1(n8911), .ip2(\cache_data[0][0] ), .op(n8166) );
  nor3_1 U8263 ( .ip1(addr_resp[7]), .ip2(addr_resp[4]), .ip3(n8158), .op(
        n12228) );
  inv_1 U8264 ( .ip(n8928), .op(n8900) );
  nand2_1 U8265 ( .ip1(n8900), .ip2(\cache_data[2][0] ), .op(n8165) );
  nor2_1 U8266 ( .ip1(n8160), .ip2(n8159), .op(n12240) );
  buf_1 U8267 ( .ip(n12240), .op(n10964) );
  nand2_1 U8268 ( .ip1(n10964), .ip2(\cache_data[5][0] ), .op(n8164) );
  nor2_1 U8269 ( .ip1(n8162), .ip2(n8161), .op(n12220) );
  buf_1 U8270 ( .ip(n12220), .op(n11971) );
  inv_1 U8271 ( .ip(n11971), .op(n11600) );
  inv_1 U8272 ( .ip(n11600), .op(n11688) );
  nand2_1 U8273 ( .ip1(n11971), .ip2(\cache_data[14][0] ), .op(n8163) );
  nand4_1 U8274 ( .ip1(n8166), .ip2(n8165), .ip3(n8164), .ip4(n8163), .op(
        n8167) );
  or4_1 U8275 ( .ip1(n8170), .ip2(n8169), .ip3(n8168), .ip4(n8167), .op(n11012) );
  nand2_1 U8276 ( .ip1(n10828), .ip2(n11012), .op(n8236) );
  nand2_1 U8277 ( .ip1(n9675), .ip2(\cache_data[5][32] ), .op(n8174) );
  nand2_1 U8278 ( .ip1(n12196), .ip2(\cache_data[10][32] ), .op(n8173) );
  nand2_1 U8279 ( .ip1(n12221), .ip2(\cache_data[15][32] ), .op(n8172) );
  nand2_1 U8280 ( .ip1(n8911), .ip2(\cache_data[0][32] ), .op(n8171) );
  nand4_1 U8281 ( .ip1(n8174), .ip2(n8173), .ip3(n8172), .ip4(n8171), .op(
        n8190) );
  nand2_1 U8282 ( .ip1(n8900), .ip2(\cache_data[2][32] ), .op(n8178) );
  nand2_1 U8283 ( .ip1(n11317), .ip2(\cache_data[3][32] ), .op(n8177) );
  nand2_1 U8284 ( .ip1(n8905), .ip2(\cache_data[6][32] ), .op(n8176) );
  nand2_1 U8285 ( .ip1(n8906), .ip2(\cache_data[4][32] ), .op(n8175) );
  nand4_1 U8286 ( .ip1(n8178), .ip2(n8177), .ip3(n8176), .ip4(n8175), .op(
        n8189) );
  nand2_1 U8287 ( .ip1(n12096), .ip2(\cache_data[11][32] ), .op(n8182) );
  nand2_1 U8288 ( .ip1(n11971), .ip2(\cache_data[14][32] ), .op(n8181) );
  nand2_1 U8289 ( .ip1(n12126), .ip2(\cache_data[9][32] ), .op(n8180) );
  nand2_1 U8290 ( .ip1(n12121), .ip2(\cache_data[8][32] ), .op(n8179) );
  nand4_1 U8291 ( .ip1(n8182), .ip2(n8181), .ip3(n8180), .ip4(n8179), .op(
        n8188) );
  nand2_1 U8292 ( .ip1(n8894), .ip2(\cache_data[1][32] ), .op(n8186) );
  nand2_1 U8293 ( .ip1(n12207), .ip2(\cache_data[12][32] ), .op(n8185) );
  nand2_1 U8294 ( .ip1(n8899), .ip2(\cache_data[13][32] ), .op(n8184) );
  nand2_1 U8295 ( .ip1(n12226), .ip2(\cache_data[7][32] ), .op(n8183) );
  nand4_1 U8296 ( .ip1(n8186), .ip2(n8185), .ip3(n8184), .ip4(n8183), .op(
        n8187) );
  nor4_1 U8297 ( .ip1(n8190), .ip2(n8189), .ip3(n8188), .ip4(n8187), .op(
        n11015) );
  nand3_1 U8298 ( .ip1(mem_data_cnt[2]), .ip2(n8211), .ip3(n11438), .op(n10870) );
  nor2_1 U8299 ( .ip1(n11015), .ip2(n10870), .op(n8213) );
  nand2_1 U8300 ( .ip1(n11971), .ip2(\cache_data[14][64] ), .op(n8194) );
  nand2_1 U8301 ( .ip1(n12126), .ip2(\cache_data[9][64] ), .op(n8193) );
  nand2_1 U8302 ( .ip1(n8900), .ip2(\cache_data[2][64] ), .op(n8192) );
  nand2_1 U8303 ( .ip1(n12207), .ip2(\cache_data[12][64] ), .op(n8191) );
  nand4_1 U8304 ( .ip1(n8194), .ip2(n8193), .ip3(n8192), .ip4(n8191), .op(
        n8210) );
  nand2_1 U8305 ( .ip1(n11317), .ip2(\cache_data[3][64] ), .op(n8198) );
  nand2_1 U8306 ( .ip1(n12196), .ip2(\cache_data[10][64] ), .op(n8197) );
  nand2_1 U8307 ( .ip1(n12221), .ip2(\cache_data[15][64] ), .op(n8196) );
  nand2_1 U8308 ( .ip1(n12240), .ip2(\cache_data[5][64] ), .op(n8195) );
  nand4_1 U8309 ( .ip1(n8198), .ip2(n8197), .ip3(n8196), .ip4(n8195), .op(
        n8209) );
  nand2_1 U8310 ( .ip1(n8894), .ip2(\cache_data[1][64] ), .op(n8202) );
  nand2_1 U8311 ( .ip1(n8905), .ip2(\cache_data[6][64] ), .op(n8201) );
  nand2_1 U8312 ( .ip1(n12121), .ip2(\cache_data[8][64] ), .op(n8200) );
  nand2_1 U8313 ( .ip1(n8906), .ip2(\cache_data[4][64] ), .op(n8199) );
  nand4_1 U8314 ( .ip1(n8202), .ip2(n8201), .ip3(n8200), .ip4(n8199), .op(
        n8208) );
  nand2_1 U8315 ( .ip1(n8911), .ip2(\cache_data[0][64] ), .op(n8206) );
  nand2_1 U8316 ( .ip1(n12226), .ip2(\cache_data[7][64] ), .op(n8205) );
  nand2_1 U8317 ( .ip1(n8899), .ip2(\cache_data[13][64] ), .op(n8204) );
  nand2_1 U8318 ( .ip1(n9669), .ip2(\cache_data[11][64] ), .op(n8203) );
  nand4_1 U8319 ( .ip1(n8206), .ip2(n8205), .ip3(n8204), .ip4(n8203), .op(
        n8207) );
  nor4_1 U8320 ( .ip1(n8210), .ip2(n8209), .ip3(n8208), .ip4(n8207), .op(
        n11013) );
  nand3_1 U8321 ( .ip1(mem_data_cnt[3]), .ip2(n8211), .ip3(n11433), .op(n10849) );
  nor2_1 U8322 ( .ip1(n11013), .ip2(n10849), .op(n8212) );
  not_ab_or_c_or_d U8323 ( .ip1(data_wr_mem[0]), .ip2(n10873), .ip3(n8213), 
        .ip4(n8212), .op(n8235) );
  nor3_1 U8324 ( .ip1(n11438), .ip2(n11433), .ip3(n10873), .op(n10894) );
  nand2_1 U8325 ( .ip1(n12226), .ip2(\cache_data[7][96] ), .op(n8217) );
  nand2_1 U8326 ( .ip1(n12121), .ip2(\cache_data[8][96] ), .op(n8216) );
  nand2_1 U8327 ( .ip1(n11971), .ip2(\cache_data[14][96] ), .op(n8215) );
  nand2_1 U8328 ( .ip1(n8906), .ip2(\cache_data[4][96] ), .op(n8214) );
  nand4_1 U8329 ( .ip1(n8217), .ip2(n8216), .ip3(n8215), .ip4(n8214), .op(
        n8233) );
  nand2_1 U8330 ( .ip1(n8894), .ip2(\cache_data[1][96] ), .op(n8221) );
  nand2_1 U8331 ( .ip1(n12096), .ip2(\cache_data[11][96] ), .op(n8220) );
  nand2_1 U8332 ( .ip1(n10975), .ip2(\cache_data[15][96] ), .op(n8219) );
  nand2_1 U8333 ( .ip1(n10964), .ip2(\cache_data[5][96] ), .op(n8218) );
  nand4_1 U8334 ( .ip1(n8221), .ip2(n8220), .ip3(n8219), .ip4(n8218), .op(
        n8232) );
  nand2_1 U8335 ( .ip1(n8900), .ip2(\cache_data[2][96] ), .op(n8225) );
  nand2_1 U8336 ( .ip1(n12196), .ip2(\cache_data[10][96] ), .op(n8224) );
  nand2_1 U8337 ( .ip1(n8905), .ip2(\cache_data[6][96] ), .op(n8223) );
  nand2_1 U8338 ( .ip1(n12207), .ip2(\cache_data[12][96] ), .op(n8222) );
  nand4_1 U8339 ( .ip1(n8225), .ip2(n8224), .ip3(n8223), .ip4(n8222), .op(
        n8231) );
  nand2_1 U8340 ( .ip1(n8911), .ip2(\cache_data[0][96] ), .op(n8229) );
  nand2_1 U8341 ( .ip1(n8899), .ip2(\cache_data[13][96] ), .op(n8228) );
  nand2_1 U8342 ( .ip1(n11317), .ip2(\cache_data[3][96] ), .op(n8227) );
  nand2_1 U8343 ( .ip1(n12126), .ip2(\cache_data[9][96] ), .op(n8226) );
  nand4_1 U8344 ( .ip1(n8229), .ip2(n8228), .ip3(n8227), .ip4(n8226), .op(
        n8230) );
  or4_1 U8345 ( .ip1(n8233), .ip2(n8232), .ip3(n8231), .ip4(n8230), .op(n11018) );
  nand2_1 U8346 ( .ip1(n10894), .ip2(n11018), .op(n8234) );
  nand3_1 U8347 ( .ip1(n8236), .ip2(n8235), .ip3(n8234), .op(n7448) );
  nand2_1 U8348 ( .ip1(n8899), .ip2(\cache_data[13][1] ), .op(n8240) );
  nand2_1 U8349 ( .ip1(n8906), .ip2(\cache_data[4][1] ), .op(n8239) );
  nand2_1 U8350 ( .ip1(n11317), .ip2(\cache_data[3][1] ), .op(n8238) );
  nand2_1 U8351 ( .ip1(n8905), .ip2(\cache_data[6][1] ), .op(n8237) );
  nand4_1 U8352 ( .ip1(n8240), .ip2(n8239), .ip3(n8238), .ip4(n8237), .op(
        n8256) );
  nand2_1 U8353 ( .ip1(n8894), .ip2(\cache_data[1][1] ), .op(n8244) );
  nand2_1 U8354 ( .ip1(n10975), .ip2(\cache_data[15][1] ), .op(n8243) );
  nand2_1 U8355 ( .ip1(n8911), .ip2(\cache_data[0][1] ), .op(n8242) );
  nand2_1 U8356 ( .ip1(n8900), .ip2(\cache_data[2][1] ), .op(n8241) );
  nand4_1 U8357 ( .ip1(n8244), .ip2(n8243), .ip3(n8242), .ip4(n8241), .op(
        n8255) );
  nand2_1 U8358 ( .ip1(n12226), .ip2(\cache_data[7][1] ), .op(n8248) );
  nand2_1 U8359 ( .ip1(n12121), .ip2(\cache_data[8][1] ), .op(n8247) );
  nand2_1 U8360 ( .ip1(n12126), .ip2(\cache_data[9][1] ), .op(n8246) );
  nand2_1 U8361 ( .ip1(n11971), .ip2(\cache_data[14][1] ), .op(n8245) );
  nand4_1 U8362 ( .ip1(n8248), .ip2(n8247), .ip3(n8246), .ip4(n8245), .op(
        n8254) );
  nand2_1 U8363 ( .ip1(n12196), .ip2(\cache_data[10][1] ), .op(n8252) );
  nand2_1 U8364 ( .ip1(n12207), .ip2(\cache_data[12][1] ), .op(n8251) );
  nand2_1 U8365 ( .ip1(n10964), .ip2(\cache_data[5][1] ), .op(n8250) );
  nand2_1 U8366 ( .ip1(n12096), .ip2(\cache_data[11][1] ), .op(n8249) );
  nand4_1 U8367 ( .ip1(n8252), .ip2(n8251), .ip3(n8250), .ip4(n8249), .op(
        n8253) );
  or4_1 U8368 ( .ip1(n8256), .ip2(n8255), .ip3(n8254), .ip4(n8253), .op(n11027) );
  nand2_1 U8369 ( .ip1(n10828), .ip2(n11027), .op(n8321) );
  nand2_1 U8370 ( .ip1(n12220), .ip2(\cache_data[14][33] ), .op(n8260) );
  nand2_1 U8371 ( .ip1(n8906), .ip2(\cache_data[4][33] ), .op(n8259) );
  nand2_1 U8372 ( .ip1(n8911), .ip2(\cache_data[0][33] ), .op(n8258) );
  nand2_1 U8373 ( .ip1(n8894), .ip2(\cache_data[1][33] ), .op(n8257) );
  nand4_1 U8374 ( .ip1(n8260), .ip2(n8259), .ip3(n8258), .ip4(n8257), .op(
        n8276) );
  nand2_1 U8375 ( .ip1(n9669), .ip2(\cache_data[11][33] ), .op(n8264) );
  nand2_1 U8376 ( .ip1(n8905), .ip2(\cache_data[6][33] ), .op(n8263) );
  nand2_1 U8377 ( .ip1(n9681), .ip2(\cache_data[15][33] ), .op(n8262) );
  nand2_1 U8378 ( .ip1(n8900), .ip2(\cache_data[2][33] ), .op(n8261) );
  nand4_1 U8379 ( .ip1(n8264), .ip2(n8263), .ip3(n8262), .ip4(n8261), .op(
        n8275) );
  nand2_1 U8380 ( .ip1(n12121), .ip2(\cache_data[8][33] ), .op(n8268) );
  nand2_1 U8381 ( .ip1(n9675), .ip2(\cache_data[5][33] ), .op(n8267) );
  nand2_1 U8382 ( .ip1(n9560), .ip2(\cache_data[12][33] ), .op(n8266) );
  nand2_1 U8383 ( .ip1(n8899), .ip2(\cache_data[13][33] ), .op(n8265) );
  nand4_1 U8384 ( .ip1(n8268), .ip2(n8267), .ip3(n8266), .ip4(n8265), .op(
        n8274) );
  nand2_1 U8385 ( .ip1(n12226), .ip2(\cache_data[7][33] ), .op(n8272) );
  nand2_1 U8386 ( .ip1(n12152), .ip2(\cache_data[9][33] ), .op(n8271) );
  nand2_1 U8387 ( .ip1(n11317), .ip2(\cache_data[3][33] ), .op(n8270) );
  nand2_1 U8388 ( .ip1(n12196), .ip2(\cache_data[10][33] ), .op(n8269) );
  nand4_1 U8389 ( .ip1(n8272), .ip2(n8271), .ip3(n8270), .ip4(n8269), .op(
        n8273) );
  nor4_1 U8390 ( .ip1(n8276), .ip2(n8275), .ip3(n8274), .ip4(n8273), .op(
        n11024) );
  nor2_1 U8391 ( .ip1(n11024), .ip2(n10870), .op(n8298) );
  nand2_1 U8392 ( .ip1(n8899), .ip2(\cache_data[13][65] ), .op(n8280) );
  nand2_1 U8393 ( .ip1(n8911), .ip2(\cache_data[0][65] ), .op(n8279) );
  nand2_1 U8394 ( .ip1(n12030), .ip2(\cache_data[12][65] ), .op(n8278) );
  nand2_1 U8395 ( .ip1(n12143), .ip2(\cache_data[7][65] ), .op(n8277) );
  nand4_1 U8396 ( .ip1(n8280), .ip2(n8279), .ip3(n8278), .ip4(n8277), .op(
        n8296) );
  nand2_1 U8397 ( .ip1(n11317), .ip2(\cache_data[3][65] ), .op(n8284) );
  nand2_1 U8398 ( .ip1(n9681), .ip2(\cache_data[15][65] ), .op(n8283) );
  nand2_1 U8399 ( .ip1(n9675), .ip2(\cache_data[5][65] ), .op(n8282) );
  nand2_1 U8400 ( .ip1(n12126), .ip2(\cache_data[9][65] ), .op(n8281) );
  nand4_1 U8401 ( .ip1(n8284), .ip2(n8283), .ip3(n8282), .ip4(n8281), .op(
        n8295) );
  nand2_1 U8402 ( .ip1(n8906), .ip2(\cache_data[4][65] ), .op(n8288) );
  nand2_1 U8403 ( .ip1(n8900), .ip2(\cache_data[2][65] ), .op(n8287) );
  nand2_1 U8404 ( .ip1(n12220), .ip2(\cache_data[14][65] ), .op(n8286) );
  nand2_1 U8405 ( .ip1(n8905), .ip2(\cache_data[6][65] ), .op(n8285) );
  nand4_1 U8406 ( .ip1(n8288), .ip2(n8287), .ip3(n8286), .ip4(n8285), .op(
        n8294) );
  nand2_1 U8407 ( .ip1(n12191), .ip2(\cache_data[8][65] ), .op(n8292) );
  nand2_1 U8408 ( .ip1(n8894), .ip2(\cache_data[1][65] ), .op(n8291) );
  nand2_1 U8409 ( .ip1(n12196), .ip2(\cache_data[10][65] ), .op(n8290) );
  nand2_1 U8410 ( .ip1(n9669), .ip2(\cache_data[11][65] ), .op(n8289) );
  nand4_1 U8411 ( .ip1(n8292), .ip2(n8291), .ip3(n8290), .ip4(n8289), .op(
        n8293) );
  nor4_1 U8412 ( .ip1(n8296), .ip2(n8295), .ip3(n8294), .ip4(n8293), .op(
        n11023) );
  nor2_1 U8413 ( .ip1(n11023), .ip2(n10849), .op(n8297) );
  not_ab_or_c_or_d U8414 ( .ip1(data_wr_mem[1]), .ip2(n10873), .ip3(n8298), 
        .ip4(n8297), .op(n8320) );
  nand2_1 U8415 ( .ip1(n8894), .ip2(\cache_data[1][97] ), .op(n8302) );
  nand2_1 U8416 ( .ip1(n12226), .ip2(\cache_data[7][97] ), .op(n8301) );
  nand2_1 U8417 ( .ip1(n12121), .ip2(\cache_data[8][97] ), .op(n8300) );
  nand2_1 U8418 ( .ip1(n8905), .ip2(\cache_data[6][97] ), .op(n8299) );
  nand4_1 U8419 ( .ip1(n8302), .ip2(n8301), .ip3(n8300), .ip4(n8299), .op(
        n8318) );
  nand2_1 U8420 ( .ip1(n11317), .ip2(\cache_data[3][97] ), .op(n8306) );
  nand2_1 U8421 ( .ip1(n8906), .ip2(\cache_data[4][97] ), .op(n8305) );
  nand2_1 U8422 ( .ip1(n12196), .ip2(\cache_data[10][97] ), .op(n8304) );
  nand2_1 U8423 ( .ip1(n11971), .ip2(\cache_data[14][97] ), .op(n8303) );
  nand4_1 U8424 ( .ip1(n8306), .ip2(n8305), .ip3(n8304), .ip4(n8303), .op(
        n8317) );
  nand2_1 U8425 ( .ip1(n8911), .ip2(\cache_data[0][97] ), .op(n8310) );
  nand2_1 U8426 ( .ip1(n12126), .ip2(\cache_data[9][97] ), .op(n8309) );
  nand2_1 U8427 ( .ip1(n12096), .ip2(\cache_data[11][97] ), .op(n8308) );
  nand2_1 U8428 ( .ip1(n12207), .ip2(\cache_data[12][97] ), .op(n8307) );
  nand4_1 U8429 ( .ip1(n8310), .ip2(n8309), .ip3(n8308), .ip4(n8307), .op(
        n8316) );
  nand2_1 U8430 ( .ip1(n8900), .ip2(\cache_data[2][97] ), .op(n8314) );
  nand2_1 U8431 ( .ip1(n10964), .ip2(\cache_data[5][97] ), .op(n8313) );
  nand2_1 U8432 ( .ip1(n10975), .ip2(\cache_data[15][97] ), .op(n8312) );
  nand2_1 U8433 ( .ip1(n8899), .ip2(\cache_data[13][97] ), .op(n8311) );
  nand4_1 U8434 ( .ip1(n8314), .ip2(n8313), .ip3(n8312), .ip4(n8311), .op(
        n8315) );
  or4_1 U8435 ( .ip1(n8318), .ip2(n8317), .ip3(n8316), .ip4(n8315), .op(n11022) );
  nand2_1 U8436 ( .ip1(n10894), .ip2(n11022), .op(n8319) );
  nand3_1 U8437 ( .ip1(n8321), .ip2(n8320), .ip3(n8319), .op(n7447) );
  nand2_1 U8438 ( .ip1(data_wr_mem[2]), .ip2(n10873), .op(n8406) );
  nand2_1 U8439 ( .ip1(n8905), .ip2(\cache_data[6][2] ), .op(n8325) );
  nand2_1 U8440 ( .ip1(n12207), .ip2(\cache_data[12][2] ), .op(n8324) );
  nand2_1 U8441 ( .ip1(n12196), .ip2(\cache_data[10][2] ), .op(n8323) );
  nand2_1 U8442 ( .ip1(n8900), .ip2(\cache_data[2][2] ), .op(n8322) );
  nand4_1 U8443 ( .ip1(n8325), .ip2(n8324), .ip3(n8323), .ip4(n8322), .op(
        n8341) );
  nand2_1 U8444 ( .ip1(n8906), .ip2(\cache_data[4][2] ), .op(n8329) );
  nand2_1 U8445 ( .ip1(n10975), .ip2(\cache_data[15][2] ), .op(n8328) );
  nand2_1 U8446 ( .ip1(n12126), .ip2(\cache_data[9][2] ), .op(n8327) );
  nand2_1 U8447 ( .ip1(n12121), .ip2(\cache_data[8][2] ), .op(n8326) );
  nand4_1 U8448 ( .ip1(n8329), .ip2(n8328), .ip3(n8327), .ip4(n8326), .op(
        n8340) );
  nand2_1 U8449 ( .ip1(n12226), .ip2(\cache_data[7][2] ), .op(n8333) );
  nand2_1 U8450 ( .ip1(n11317), .ip2(\cache_data[3][2] ), .op(n8332) );
  nand2_1 U8451 ( .ip1(n12096), .ip2(\cache_data[11][2] ), .op(n8331) );
  nand2_1 U8452 ( .ip1(n8894), .ip2(\cache_data[1][2] ), .op(n8330) );
  nand4_1 U8453 ( .ip1(n8333), .ip2(n8332), .ip3(n8331), .ip4(n8330), .op(
        n8339) );
  nand2_1 U8454 ( .ip1(n8911), .ip2(\cache_data[0][2] ), .op(n8337) );
  nand2_1 U8455 ( .ip1(n8899), .ip2(\cache_data[13][2] ), .op(n8336) );
  nand2_1 U8456 ( .ip1(n11971), .ip2(\cache_data[14][2] ), .op(n8335) );
  nand2_1 U8457 ( .ip1(n10964), .ip2(\cache_data[5][2] ), .op(n8334) );
  nand4_1 U8458 ( .ip1(n8337), .ip2(n8336), .ip3(n8335), .ip4(n8334), .op(
        n8338) );
  or4_1 U8459 ( .ip1(n8341), .ip2(n8340), .ip3(n8339), .ip4(n8338), .op(n11031) );
  nand2_1 U8460 ( .ip1(n12126), .ip2(\cache_data[9][66] ), .op(n8345) );
  nand2_1 U8461 ( .ip1(n12196), .ip2(\cache_data[10][66] ), .op(n8344) );
  nand2_1 U8462 ( .ip1(n12226), .ip2(\cache_data[7][66] ), .op(n8343) );
  nand2_1 U8463 ( .ip1(n8911), .ip2(\cache_data[0][66] ), .op(n8342) );
  nand4_1 U8464 ( .ip1(n8345), .ip2(n8344), .ip3(n8343), .ip4(n8342), .op(
        n8361) );
  nand2_1 U8465 ( .ip1(n9681), .ip2(\cache_data[15][66] ), .op(n8349) );
  nand2_1 U8466 ( .ip1(n11317), .ip2(\cache_data[3][66] ), .op(n8348) );
  nand2_1 U8467 ( .ip1(n12191), .ip2(\cache_data[8][66] ), .op(n8347) );
  nand2_1 U8468 ( .ip1(n12207), .ip2(\cache_data[12][66] ), .op(n8346) );
  nand4_1 U8469 ( .ip1(n8349), .ip2(n8348), .ip3(n8347), .ip4(n8346), .op(
        n8360) );
  nand2_1 U8470 ( .ip1(n8905), .ip2(\cache_data[6][66] ), .op(n8353) );
  nand2_1 U8471 ( .ip1(n11971), .ip2(\cache_data[14][66] ), .op(n8352) );
  nand2_1 U8472 ( .ip1(n8906), .ip2(\cache_data[4][66] ), .op(n8351) );
  nand2_1 U8473 ( .ip1(n8894), .ip2(\cache_data[1][66] ), .op(n8350) );
  nand4_1 U8474 ( .ip1(n8353), .ip2(n8352), .ip3(n8351), .ip4(n8350), .op(
        n8359) );
  nand2_1 U8475 ( .ip1(n9669), .ip2(\cache_data[11][66] ), .op(n8357) );
  nand2_1 U8476 ( .ip1(n9675), .ip2(\cache_data[5][66] ), .op(n8356) );
  nand2_1 U8477 ( .ip1(n8899), .ip2(\cache_data[13][66] ), .op(n8355) );
  nand2_1 U8478 ( .ip1(n8900), .ip2(\cache_data[2][66] ), .op(n8354) );
  nand4_1 U8479 ( .ip1(n8357), .ip2(n8356), .ip3(n8355), .ip4(n8354), .op(
        n8358) );
  nor4_1 U8480 ( .ip1(n8361), .ip2(n8360), .ip3(n8359), .ip4(n8358), .op(
        n11032) );
  nor2_1 U8481 ( .ip1(n11032), .ip2(n10849), .op(n8383) );
  nand2_1 U8482 ( .ip1(n8894), .ip2(\cache_data[1][34] ), .op(n8365) );
  nand2_1 U8483 ( .ip1(n11317), .ip2(\cache_data[3][34] ), .op(n8364) );
  nand2_1 U8484 ( .ip1(n8899), .ip2(\cache_data[13][34] ), .op(n8363) );
  nand2_1 U8485 ( .ip1(n9681), .ip2(\cache_data[15][34] ), .op(n8362) );
  nand4_1 U8486 ( .ip1(n8365), .ip2(n8364), .ip3(n8363), .ip4(n8362), .op(
        n8381) );
  nand2_1 U8487 ( .ip1(n12096), .ip2(\cache_data[11][34] ), .op(n8369) );
  nand2_1 U8488 ( .ip1(n8900), .ip2(\cache_data[2][34] ), .op(n8368) );
  nand2_1 U8489 ( .ip1(n12207), .ip2(\cache_data[12][34] ), .op(n8367) );
  nand2_1 U8490 ( .ip1(n8905), .ip2(\cache_data[6][34] ), .op(n8366) );
  nand4_1 U8491 ( .ip1(n8369), .ip2(n8368), .ip3(n8367), .ip4(n8366), .op(
        n8380) );
  nand2_1 U8492 ( .ip1(n10964), .ip2(\cache_data[5][34] ), .op(n8373) );
  nand2_1 U8493 ( .ip1(n12196), .ip2(\cache_data[10][34] ), .op(n8372) );
  nand2_1 U8494 ( .ip1(n11971), .ip2(\cache_data[14][34] ), .op(n8371) );
  nand2_1 U8495 ( .ip1(n12226), .ip2(\cache_data[7][34] ), .op(n8370) );
  nand4_1 U8496 ( .ip1(n8373), .ip2(n8372), .ip3(n8371), .ip4(n8370), .op(
        n8379) );
  nand2_1 U8497 ( .ip1(n12121), .ip2(\cache_data[8][34] ), .op(n8377) );
  nand2_1 U8498 ( .ip1(n8906), .ip2(\cache_data[4][34] ), .op(n8376) );
  nand2_1 U8499 ( .ip1(n8911), .ip2(\cache_data[0][34] ), .op(n8375) );
  nand2_1 U8500 ( .ip1(n9682), .ip2(\cache_data[9][34] ), .op(n8374) );
  nand4_1 U8501 ( .ip1(n8377), .ip2(n8376), .ip3(n8375), .ip4(n8374), .op(
        n8378) );
  nor4_1 U8502 ( .ip1(n8381), .ip2(n8380), .ip3(n8379), .ip4(n8378), .op(
        n11033) );
  nor2_1 U8503 ( .ip1(n11033), .ip2(n10870), .op(n8382) );
  not_ab_or_c_or_d U8504 ( .ip1(n10828), .ip2(n11031), .ip3(n8383), .ip4(n8382), .op(n8405) );
  nand2_1 U8505 ( .ip1(n12096), .ip2(\cache_data[11][98] ), .op(n8387) );
  nand2_1 U8506 ( .ip1(n12196), .ip2(\cache_data[10][98] ), .op(n8386) );
  nand2_1 U8507 ( .ip1(n8911), .ip2(\cache_data[0][98] ), .op(n8385) );
  nand2_1 U8508 ( .ip1(n12121), .ip2(\cache_data[8][98] ), .op(n8384) );
  nand4_1 U8509 ( .ip1(n8387), .ip2(n8386), .ip3(n8385), .ip4(n8384), .op(
        n8403) );
  nand2_1 U8510 ( .ip1(n8900), .ip2(\cache_data[2][98] ), .op(n8391) );
  nand2_1 U8511 ( .ip1(n12226), .ip2(\cache_data[7][98] ), .op(n8390) );
  nand2_1 U8512 ( .ip1(n10975), .ip2(\cache_data[15][98] ), .op(n8389) );
  nand2_1 U8513 ( .ip1(n12207), .ip2(\cache_data[12][98] ), .op(n8388) );
  nand4_1 U8514 ( .ip1(n8391), .ip2(n8390), .ip3(n8389), .ip4(n8388), .op(
        n8402) );
  nand2_1 U8515 ( .ip1(n8906), .ip2(\cache_data[4][98] ), .op(n8395) );
  nand2_1 U8516 ( .ip1(n12126), .ip2(\cache_data[9][98] ), .op(n8394) );
  nand2_1 U8517 ( .ip1(n11317), .ip2(\cache_data[3][98] ), .op(n8393) );
  nand2_1 U8518 ( .ip1(n11971), .ip2(\cache_data[14][98] ), .op(n8392) );
  nand4_1 U8519 ( .ip1(n8395), .ip2(n8394), .ip3(n8393), .ip4(n8392), .op(
        n8401) );
  nand2_1 U8520 ( .ip1(n10964), .ip2(\cache_data[5][98] ), .op(n8399) );
  nand2_1 U8521 ( .ip1(n8899), .ip2(\cache_data[13][98] ), .op(n8398) );
  nand2_1 U8522 ( .ip1(n8905), .ip2(\cache_data[6][98] ), .op(n8397) );
  nand2_1 U8523 ( .ip1(n8894), .ip2(\cache_data[1][98] ), .op(n8396) );
  nand4_1 U8524 ( .ip1(n8399), .ip2(n8398), .ip3(n8397), .ip4(n8396), .op(
        n8400) );
  or4_1 U8525 ( .ip1(n8403), .ip2(n8402), .ip3(n8401), .ip4(n8400), .op(n11036) );
  nand2_1 U8526 ( .ip1(n10894), .ip2(n11036), .op(n8404) );
  nand3_1 U8527 ( .ip1(n8406), .ip2(n8405), .ip3(n8404), .op(n7446) );
  nand2_1 U8528 ( .ip1(n8894), .ip2(\cache_data[1][3] ), .op(n8410) );
  nand2_1 U8529 ( .ip1(n12126), .ip2(\cache_data[9][3] ), .op(n8409) );
  nand2_1 U8530 ( .ip1(n11317), .ip2(\cache_data[3][3] ), .op(n8408) );
  nand2_1 U8531 ( .ip1(n12220), .ip2(\cache_data[14][3] ), .op(n8407) );
  nand4_1 U8532 ( .ip1(n8410), .ip2(n8409), .ip3(n8408), .ip4(n8407), .op(
        n8426) );
  nand2_1 U8533 ( .ip1(n12226), .ip2(\cache_data[7][3] ), .op(n8414) );
  nand2_1 U8534 ( .ip1(n8899), .ip2(\cache_data[13][3] ), .op(n8413) );
  nand2_1 U8535 ( .ip1(n8906), .ip2(\cache_data[4][3] ), .op(n8412) );
  nand2_1 U8536 ( .ip1(n10975), .ip2(\cache_data[15][3] ), .op(n8411) );
  nand4_1 U8537 ( .ip1(n8414), .ip2(n8413), .ip3(n8412), .ip4(n8411), .op(
        n8425) );
  nand2_1 U8538 ( .ip1(n10964), .ip2(\cache_data[5][3] ), .op(n8418) );
  nand2_1 U8539 ( .ip1(n12207), .ip2(\cache_data[12][3] ), .op(n8417) );
  nand2_1 U8540 ( .ip1(n8905), .ip2(\cache_data[6][3] ), .op(n8416) );
  nand2_1 U8541 ( .ip1(n12096), .ip2(\cache_data[11][3] ), .op(n8415) );
  nand4_1 U8542 ( .ip1(n8418), .ip2(n8417), .ip3(n8416), .ip4(n8415), .op(
        n8424) );
  nand2_1 U8543 ( .ip1(n8911), .ip2(\cache_data[0][3] ), .op(n8422) );
  nand2_1 U8544 ( .ip1(n8900), .ip2(\cache_data[2][3] ), .op(n8421) );
  nand2_1 U8545 ( .ip1(n12235), .ip2(\cache_data[10][3] ), .op(n8420) );
  nand2_1 U8546 ( .ip1(n12121), .ip2(\cache_data[8][3] ), .op(n8419) );
  nand4_1 U8547 ( .ip1(n8422), .ip2(n8421), .ip3(n8420), .ip4(n8419), .op(
        n8423) );
  or4_1 U8548 ( .ip1(n8426), .ip2(n8425), .ip3(n8424), .ip4(n8423), .op(n11040) );
  nand2_1 U8549 ( .ip1(n10828), .ip2(n11040), .op(n8491) );
  nand2_1 U8550 ( .ip1(n8900), .ip2(\cache_data[2][67] ), .op(n8430) );
  nand2_1 U8551 ( .ip1(n12121), .ip2(\cache_data[8][67] ), .op(n8429) );
  nand2_1 U8552 ( .ip1(n12226), .ip2(\cache_data[7][67] ), .op(n8428) );
  nand2_1 U8553 ( .ip1(n12220), .ip2(\cache_data[14][67] ), .op(n8427) );
  nand4_1 U8554 ( .ip1(n8430), .ip2(n8429), .ip3(n8428), .ip4(n8427), .op(
        n8446) );
  nand2_1 U8555 ( .ip1(n12196), .ip2(\cache_data[10][67] ), .op(n8434) );
  nand2_1 U8556 ( .ip1(n11317), .ip2(\cache_data[3][67] ), .op(n8433) );
  nand2_1 U8557 ( .ip1(n8899), .ip2(\cache_data[13][67] ), .op(n8432) );
  nand2_1 U8558 ( .ip1(n8894), .ip2(\cache_data[1][67] ), .op(n8431) );
  nand4_1 U8559 ( .ip1(n8434), .ip2(n8433), .ip3(n8432), .ip4(n8431), .op(
        n8445) );
  nand2_1 U8560 ( .ip1(n8906), .ip2(\cache_data[4][67] ), .op(n8438) );
  nand2_1 U8561 ( .ip1(n8911), .ip2(\cache_data[0][67] ), .op(n8437) );
  nand2_1 U8562 ( .ip1(n9681), .ip2(\cache_data[15][67] ), .op(n8436) );
  nand2_1 U8563 ( .ip1(n9669), .ip2(\cache_data[11][67] ), .op(n8435) );
  nand4_1 U8564 ( .ip1(n8438), .ip2(n8437), .ip3(n8436), .ip4(n8435), .op(
        n8444) );
  nand2_1 U8565 ( .ip1(n12241), .ip2(\cache_data[9][67] ), .op(n8442) );
  nand2_1 U8566 ( .ip1(n12227), .ip2(\cache_data[12][67] ), .op(n8441) );
  nand2_1 U8567 ( .ip1(n9675), .ip2(\cache_data[5][67] ), .op(n8440) );
  nand2_1 U8568 ( .ip1(n8905), .ip2(\cache_data[6][67] ), .op(n8439) );
  nand4_1 U8569 ( .ip1(n8442), .ip2(n8441), .ip3(n8440), .ip4(n8439), .op(
        n8443) );
  nor4_1 U8570 ( .ip1(n8446), .ip2(n8445), .ip3(n8444), .ip4(n8443), .op(
        n11042) );
  nor2_1 U8571 ( .ip1(n11042), .ip2(n10849), .op(n8468) );
  nand2_1 U8572 ( .ip1(n12235), .ip2(\cache_data[10][35] ), .op(n8450) );
  nand2_1 U8573 ( .ip1(n9669), .ip2(\cache_data[11][35] ), .op(n8449) );
  nand2_1 U8574 ( .ip1(n8911), .ip2(\cache_data[0][35] ), .op(n8448) );
  nand2_1 U8575 ( .ip1(n12226), .ip2(\cache_data[7][35] ), .op(n8447) );
  nand4_1 U8576 ( .ip1(n8450), .ip2(n8449), .ip3(n8448), .ip4(n8447), .op(
        n8466) );
  nand2_1 U8577 ( .ip1(n8899), .ip2(\cache_data[13][35] ), .op(n8454) );
  nand2_1 U8578 ( .ip1(n10975), .ip2(\cache_data[15][35] ), .op(n8453) );
  nand2_1 U8579 ( .ip1(n11317), .ip2(\cache_data[3][35] ), .op(n8452) );
  nand2_1 U8580 ( .ip1(n8906), .ip2(\cache_data[4][35] ), .op(n8451) );
  nand4_1 U8581 ( .ip1(n8454), .ip2(n8453), .ip3(n8452), .ip4(n8451), .op(
        n8465) );
  nand2_1 U8582 ( .ip1(n8905), .ip2(\cache_data[6][35] ), .op(n8458) );
  nand2_1 U8583 ( .ip1(n9675), .ip2(\cache_data[5][35] ), .op(n8457) );
  nand2_1 U8584 ( .ip1(n12220), .ip2(\cache_data[14][35] ), .op(n8456) );
  nand2_1 U8585 ( .ip1(n12120), .ip2(\cache_data[1][35] ), .op(n8455) );
  nand4_1 U8586 ( .ip1(n8458), .ip2(n8457), .ip3(n8456), .ip4(n8455), .op(
        n8464) );
  nand2_1 U8587 ( .ip1(n12121), .ip2(\cache_data[8][35] ), .op(n8462) );
  nand2_1 U8588 ( .ip1(n9560), .ip2(\cache_data[12][35] ), .op(n8461) );
  nand2_1 U8589 ( .ip1(n8900), .ip2(\cache_data[2][35] ), .op(n8460) );
  nand2_1 U8590 ( .ip1(n12241), .ip2(\cache_data[9][35] ), .op(n8459) );
  nand4_1 U8591 ( .ip1(n8462), .ip2(n8461), .ip3(n8460), .ip4(n8459), .op(
        n8463) );
  nor4_1 U8592 ( .ip1(n8466), .ip2(n8465), .ip3(n8464), .ip4(n8463), .op(
        n11041) );
  nor2_1 U8593 ( .ip1(n11041), .ip2(n10870), .op(n8467) );
  not_ab_or_c_or_d U8594 ( .ip1(data_wr_mem[3]), .ip2(n10873), .ip3(n8468), 
        .ip4(n8467), .op(n8490) );
  nand2_1 U8595 ( .ip1(n12235), .ip2(\cache_data[10][99] ), .op(n8472) );
  nand2_1 U8596 ( .ip1(n12096), .ip2(\cache_data[11][99] ), .op(n8471) );
  nand2_1 U8597 ( .ip1(n8911), .ip2(\cache_data[0][99] ), .op(n8470) );
  nand2_1 U8598 ( .ip1(n12121), .ip2(\cache_data[8][99] ), .op(n8469) );
  nand4_1 U8599 ( .ip1(n8472), .ip2(n8471), .ip3(n8470), .ip4(n8469), .op(
        n8488) );
  nand2_1 U8600 ( .ip1(n12220), .ip2(\cache_data[14][99] ), .op(n8476) );
  nand2_1 U8601 ( .ip1(n12207), .ip2(\cache_data[12][99] ), .op(n8475) );
  nand2_1 U8602 ( .ip1(n10975), .ip2(\cache_data[15][99] ), .op(n8474) );
  nand2_1 U8603 ( .ip1(n11317), .ip2(\cache_data[3][99] ), .op(n8473) );
  nand4_1 U8604 ( .ip1(n8476), .ip2(n8475), .ip3(n8474), .ip4(n8473), .op(
        n8487) );
  nand2_1 U8605 ( .ip1(n8905), .ip2(\cache_data[6][99] ), .op(n8480) );
  nand2_1 U8606 ( .ip1(n8899), .ip2(\cache_data[13][99] ), .op(n8479) );
  nand2_1 U8607 ( .ip1(n8900), .ip2(\cache_data[2][99] ), .op(n8478) );
  nand2_1 U8608 ( .ip1(n8906), .ip2(\cache_data[4][99] ), .op(n8477) );
  nand4_1 U8609 ( .ip1(n8480), .ip2(n8479), .ip3(n8478), .ip4(n8477), .op(
        n8486) );
  nand2_1 U8610 ( .ip1(n8894), .ip2(\cache_data[1][99] ), .op(n8484) );
  nand2_1 U8611 ( .ip1(n12241), .ip2(\cache_data[9][99] ), .op(n8483) );
  nand2_1 U8612 ( .ip1(n10964), .ip2(\cache_data[5][99] ), .op(n8482) );
  nand2_1 U8613 ( .ip1(n12226), .ip2(\cache_data[7][99] ), .op(n8481) );
  nand4_1 U8614 ( .ip1(n8484), .ip2(n8483), .ip3(n8482), .ip4(n8481), .op(
        n8485) );
  or4_1 U8615 ( .ip1(n8488), .ip2(n8487), .ip3(n8486), .ip4(n8485), .op(n11045) );
  nand2_1 U8616 ( .ip1(n10894), .ip2(n11045), .op(n8489) );
  nand3_1 U8617 ( .ip1(n8491), .ip2(n8490), .ip3(n8489), .op(n7445) );
  nand2_1 U8618 ( .ip1(data_wr_mem[4]), .ip2(n10873), .op(n8576) );
  nand2_1 U8619 ( .ip1(n12207), .ip2(\cache_data[12][100] ), .op(n8495) );
  nand2_1 U8620 ( .ip1(n10975), .ip2(\cache_data[15][100] ), .op(n8494) );
  nand2_1 U8621 ( .ip1(n8899), .ip2(\cache_data[13][100] ), .op(n8493) );
  nand2_1 U8622 ( .ip1(n10964), .ip2(\cache_data[5][100] ), .op(n8492) );
  nand4_1 U8623 ( .ip1(n8495), .ip2(n8494), .ip3(n8493), .ip4(n8492), .op(
        n8511) );
  nand2_1 U8624 ( .ip1(n8905), .ip2(\cache_data[6][100] ), .op(n8499) );
  nand2_1 U8625 ( .ip1(n8900), .ip2(\cache_data[2][100] ), .op(n8498) );
  nand2_1 U8626 ( .ip1(n12241), .ip2(\cache_data[9][100] ), .op(n8497) );
  nand2_1 U8627 ( .ip1(n12096), .ip2(\cache_data[11][100] ), .op(n8496) );
  nand4_1 U8628 ( .ip1(n8499), .ip2(n8498), .ip3(n8497), .ip4(n8496), .op(
        n8510) );
  nand2_1 U8629 ( .ip1(n12121), .ip2(\cache_data[8][100] ), .op(n8503) );
  nand2_1 U8630 ( .ip1(n12220), .ip2(\cache_data[14][100] ), .op(n8502) );
  nand2_1 U8631 ( .ip1(n8911), .ip2(\cache_data[0][100] ), .op(n8501) );
  nand2_1 U8632 ( .ip1(n12235), .ip2(\cache_data[10][100] ), .op(n8500) );
  nand4_1 U8633 ( .ip1(n8503), .ip2(n8502), .ip3(n8501), .ip4(n8500), .op(
        n8509) );
  nand2_1 U8634 ( .ip1(n12226), .ip2(\cache_data[7][100] ), .op(n8507) );
  nand2_1 U8635 ( .ip1(n8906), .ip2(\cache_data[4][100] ), .op(n8506) );
  nand2_1 U8636 ( .ip1(n12120), .ip2(\cache_data[1][100] ), .op(n8505) );
  nand2_1 U8637 ( .ip1(n11317), .ip2(\cache_data[3][100] ), .op(n8504) );
  nand4_1 U8638 ( .ip1(n8507), .ip2(n8506), .ip3(n8505), .ip4(n8504), .op(
        n8508) );
  or4_1 U8639 ( .ip1(n8511), .ip2(n8510), .ip3(n8509), .ip4(n8508), .op(n11049) );
  nand2_1 U8640 ( .ip1(n8905), .ip2(\cache_data[6][36] ), .op(n8515) );
  nand2_1 U8641 ( .ip1(n12207), .ip2(\cache_data[12][36] ), .op(n8514) );
  nand2_1 U8642 ( .ip1(n9675), .ip2(\cache_data[5][36] ), .op(n8513) );
  nand2_1 U8643 ( .ip1(n12241), .ip2(\cache_data[9][36] ), .op(n8512) );
  nand4_1 U8644 ( .ip1(n8515), .ip2(n8514), .ip3(n8513), .ip4(n8512), .op(
        n8531) );
  nand2_1 U8645 ( .ip1(n8911), .ip2(\cache_data[0][36] ), .op(n8519) );
  nand2_1 U8646 ( .ip1(n8906), .ip2(\cache_data[4][36] ), .op(n8518) );
  nand2_1 U8647 ( .ip1(n8899), .ip2(\cache_data[13][36] ), .op(n8517) );
  nand2_1 U8648 ( .ip1(n11317), .ip2(\cache_data[3][36] ), .op(n8516) );
  nand4_1 U8649 ( .ip1(n8519), .ip2(n8518), .ip3(n8517), .ip4(n8516), .op(
        n8530) );
  nand2_1 U8650 ( .ip1(n12170), .ip2(\cache_data[11][36] ), .op(n8523) );
  nand2_1 U8651 ( .ip1(n12220), .ip2(\cache_data[14][36] ), .op(n8522) );
  nand2_1 U8652 ( .ip1(n8900), .ip2(\cache_data[2][36] ), .op(n8521) );
  nand2_1 U8653 ( .ip1(n8894), .ip2(\cache_data[1][36] ), .op(n8520) );
  nand4_1 U8654 ( .ip1(n8523), .ip2(n8522), .ip3(n8521), .ip4(n8520), .op(
        n8529) );
  nand2_1 U8655 ( .ip1(n9681), .ip2(\cache_data[15][36] ), .op(n8527) );
  nand2_1 U8656 ( .ip1(n12196), .ip2(\cache_data[10][36] ), .op(n8526) );
  nand2_1 U8657 ( .ip1(n12121), .ip2(\cache_data[8][36] ), .op(n8525) );
  nand2_1 U8658 ( .ip1(n12226), .ip2(\cache_data[7][36] ), .op(n8524) );
  nand4_1 U8659 ( .ip1(n8527), .ip2(n8526), .ip3(n8525), .ip4(n8524), .op(
        n8528) );
  nor4_1 U8660 ( .ip1(n8531), .ip2(n8530), .ip3(n8529), .ip4(n8528), .op(
        n11050) );
  nor2_1 U8661 ( .ip1(n11050), .ip2(n10870), .op(n8553) );
  nand2_1 U8662 ( .ip1(n11317), .ip2(\cache_data[3][68] ), .op(n8535) );
  nand2_1 U8663 ( .ip1(n8899), .ip2(\cache_data[13][68] ), .op(n8534) );
  nand2_1 U8664 ( .ip1(n12241), .ip2(\cache_data[9][68] ), .op(n8533) );
  nand2_1 U8665 ( .ip1(n11927), .ip2(\cache_data[11][68] ), .op(n8532) );
  nand4_1 U8666 ( .ip1(n8535), .ip2(n8534), .ip3(n8533), .ip4(n8532), .op(
        n8551) );
  nand2_1 U8667 ( .ip1(n9681), .ip2(\cache_data[15][68] ), .op(n8539) );
  nand2_1 U8668 ( .ip1(n12121), .ip2(\cache_data[8][68] ), .op(n8538) );
  nand2_1 U8669 ( .ip1(n12226), .ip2(\cache_data[7][68] ), .op(n8537) );
  nand2_1 U8670 ( .ip1(n8911), .ip2(\cache_data[0][68] ), .op(n8536) );
  nand4_1 U8671 ( .ip1(n8539), .ip2(n8538), .ip3(n8537), .ip4(n8536), .op(
        n8550) );
  nand2_1 U8672 ( .ip1(n9675), .ip2(\cache_data[5][68] ), .op(n8543) );
  nand2_1 U8673 ( .ip1(n8905), .ip2(\cache_data[6][68] ), .op(n8542) );
  nand2_1 U8674 ( .ip1(n12207), .ip2(\cache_data[12][68] ), .op(n8541) );
  nand2_1 U8675 ( .ip1(n11971), .ip2(\cache_data[14][68] ), .op(n8540) );
  nand4_1 U8676 ( .ip1(n8543), .ip2(n8542), .ip3(n8541), .ip4(n8540), .op(
        n8549) );
  nand2_1 U8677 ( .ip1(n12235), .ip2(\cache_data[10][68] ), .op(n8547) );
  nand2_1 U8678 ( .ip1(n8906), .ip2(\cache_data[4][68] ), .op(n8546) );
  nand2_1 U8679 ( .ip1(n8900), .ip2(\cache_data[2][68] ), .op(n8545) );
  nand2_1 U8680 ( .ip1(n8894), .ip2(\cache_data[1][68] ), .op(n8544) );
  nand4_1 U8681 ( .ip1(n8547), .ip2(n8546), .ip3(n8545), .ip4(n8544), .op(
        n8548) );
  nor4_1 U8682 ( .ip1(n8551), .ip2(n8550), .ip3(n8549), .ip4(n8548), .op(
        n11051) );
  nor2_1 U8683 ( .ip1(n11051), .ip2(n10849), .op(n8552) );
  not_ab_or_c_or_d U8684 ( .ip1(n10894), .ip2(n11049), .ip3(n8553), .ip4(n8552), .op(n8575) );
  nand2_1 U8685 ( .ip1(n12235), .ip2(\cache_data[10][4] ), .op(n8557) );
  nand2_1 U8686 ( .ip1(n11317), .ip2(\cache_data[3][4] ), .op(n8556) );
  nand2_1 U8687 ( .ip1(n12220), .ip2(\cache_data[14][4] ), .op(n8555) );
  nand2_1 U8688 ( .ip1(n8905), .ip2(\cache_data[6][4] ), .op(n8554) );
  nand4_1 U8689 ( .ip1(n8557), .ip2(n8556), .ip3(n8555), .ip4(n8554), .op(
        n8573) );
  nand2_1 U8690 ( .ip1(n8894), .ip2(\cache_data[1][4] ), .op(n8561) );
  nand2_1 U8691 ( .ip1(n10975), .ip2(\cache_data[15][4] ), .op(n8560) );
  nand2_1 U8692 ( .ip1(n12096), .ip2(\cache_data[11][4] ), .op(n8559) );
  nand2_1 U8693 ( .ip1(n8911), .ip2(\cache_data[0][4] ), .op(n8558) );
  nand4_1 U8694 ( .ip1(n8561), .ip2(n8560), .ip3(n8559), .ip4(n8558), .op(
        n8572) );
  nand2_1 U8695 ( .ip1(n12226), .ip2(\cache_data[7][4] ), .op(n8565) );
  nand2_1 U8696 ( .ip1(n8899), .ip2(\cache_data[13][4] ), .op(n8564) );
  nand2_1 U8697 ( .ip1(n10964), .ip2(\cache_data[5][4] ), .op(n8563) );
  nand2_1 U8698 ( .ip1(n12126), .ip2(\cache_data[9][4] ), .op(n8562) );
  nand4_1 U8699 ( .ip1(n8565), .ip2(n8564), .ip3(n8563), .ip4(n8562), .op(
        n8571) );
  nand2_1 U8700 ( .ip1(n8906), .ip2(\cache_data[4][4] ), .op(n8569) );
  nand2_1 U8701 ( .ip1(n12207), .ip2(\cache_data[12][4] ), .op(n8568) );
  nand2_1 U8702 ( .ip1(n8900), .ip2(\cache_data[2][4] ), .op(n8567) );
  nand2_1 U8703 ( .ip1(n12121), .ip2(\cache_data[8][4] ), .op(n8566) );
  nand4_1 U8704 ( .ip1(n8569), .ip2(n8568), .ip3(n8567), .ip4(n8566), .op(
        n8570) );
  or4_1 U8705 ( .ip1(n8573), .ip2(n8572), .ip3(n8571), .ip4(n8570), .op(n11054) );
  nand2_1 U8706 ( .ip1(n10828), .ip2(n11054), .op(n8574) );
  nand3_1 U8707 ( .ip1(n8576), .ip2(n8575), .ip3(n8574), .op(n7444) );
  nand2_1 U8708 ( .ip1(data_wr_mem[5]), .ip2(n10873), .op(n8661) );
  nand2_1 U8709 ( .ip1(n8899), .ip2(\cache_data[13][101] ), .op(n8580) );
  nand2_1 U8710 ( .ip1(n8911), .ip2(\cache_data[0][101] ), .op(n8579) );
  nand2_1 U8711 ( .ip1(n8906), .ip2(\cache_data[4][101] ), .op(n8578) );
  nand2_1 U8712 ( .ip1(n8900), .ip2(\cache_data[2][101] ), .op(n8577) );
  nand4_1 U8713 ( .ip1(n8580), .ip2(n8579), .ip3(n8578), .ip4(n8577), .op(
        n8596) );
  nand2_1 U8714 ( .ip1(n12207), .ip2(\cache_data[12][101] ), .op(n8584) );
  nand2_1 U8715 ( .ip1(n11317), .ip2(\cache_data[3][101] ), .op(n8583) );
  nand2_1 U8716 ( .ip1(n12096), .ip2(\cache_data[11][101] ), .op(n8582) );
  nand2_1 U8717 ( .ip1(n12120), .ip2(\cache_data[1][101] ), .op(n8581) );
  nand4_1 U8718 ( .ip1(n8584), .ip2(n8583), .ip3(n8582), .ip4(n8581), .op(
        n8595) );
  nand2_1 U8719 ( .ip1(n12121), .ip2(\cache_data[8][101] ), .op(n8588) );
  nand2_1 U8720 ( .ip1(n10964), .ip2(\cache_data[5][101] ), .op(n8587) );
  nand2_1 U8721 ( .ip1(n10975), .ip2(\cache_data[15][101] ), .op(n8586) );
  nand2_1 U8722 ( .ip1(n12235), .ip2(\cache_data[10][101] ), .op(n8585) );
  nand4_1 U8723 ( .ip1(n8588), .ip2(n8587), .ip3(n8586), .ip4(n8585), .op(
        n8594) );
  nand2_1 U8724 ( .ip1(n12241), .ip2(\cache_data[9][101] ), .op(n8592) );
  nand2_1 U8725 ( .ip1(n12226), .ip2(\cache_data[7][101] ), .op(n8591) );
  nand2_1 U8726 ( .ip1(n8905), .ip2(\cache_data[6][101] ), .op(n8590) );
  nand2_1 U8727 ( .ip1(n12220), .ip2(\cache_data[14][101] ), .op(n8589) );
  nand4_1 U8728 ( .ip1(n8592), .ip2(n8591), .ip3(n8590), .ip4(n8589), .op(
        n8593) );
  or4_1 U8729 ( .ip1(n8596), .ip2(n8595), .ip3(n8594), .ip4(n8593), .op(n11058) );
  nand2_1 U8730 ( .ip1(n8906), .ip2(\cache_data[4][37] ), .op(n8600) );
  nand2_1 U8731 ( .ip1(n8899), .ip2(\cache_data[13][37] ), .op(n8599) );
  nand2_1 U8732 ( .ip1(n8911), .ip2(\cache_data[0][37] ), .op(n8598) );
  nand2_1 U8733 ( .ip1(n12202), .ip2(\cache_data[7][37] ), .op(n8597) );
  nand4_1 U8734 ( .ip1(n8600), .ip2(n8599), .ip3(n8598), .ip4(n8597), .op(
        n8616) );
  nand2_1 U8735 ( .ip1(n12207), .ip2(\cache_data[12][37] ), .op(n8604) );
  nand2_1 U8736 ( .ip1(n8894), .ip2(\cache_data[1][37] ), .op(n8603) );
  nand2_1 U8737 ( .ip1(n11317), .ip2(\cache_data[3][37] ), .op(n8602) );
  nand2_1 U8738 ( .ip1(n9675), .ip2(\cache_data[5][37] ), .op(n8601) );
  nand4_1 U8739 ( .ip1(n8604), .ip2(n8603), .ip3(n8602), .ip4(n8601), .op(
        n8615) );
  nand2_1 U8740 ( .ip1(n12121), .ip2(\cache_data[8][37] ), .op(n8608) );
  nand2_1 U8741 ( .ip1(n8905), .ip2(\cache_data[6][37] ), .op(n8607) );
  nand2_1 U8742 ( .ip1(n9669), .ip2(\cache_data[11][37] ), .op(n8606) );
  nand2_1 U8743 ( .ip1(n8900), .ip2(\cache_data[2][37] ), .op(n8605) );
  nand4_1 U8744 ( .ip1(n8608), .ip2(n8607), .ip3(n8606), .ip4(n8605), .op(
        n8614) );
  nand2_1 U8745 ( .ip1(n12235), .ip2(\cache_data[10][37] ), .op(n8612) );
  nand2_1 U8746 ( .ip1(n12241), .ip2(\cache_data[9][37] ), .op(n8611) );
  nand2_1 U8747 ( .ip1(n11971), .ip2(\cache_data[14][37] ), .op(n8610) );
  nand2_1 U8748 ( .ip1(n9681), .ip2(\cache_data[15][37] ), .op(n8609) );
  nand4_1 U8749 ( .ip1(n8612), .ip2(n8611), .ip3(n8610), .ip4(n8609), .op(
        n8613) );
  nor4_1 U8750 ( .ip1(n8616), .ip2(n8615), .ip3(n8614), .ip4(n8613), .op(
        n11060) );
  nor2_1 U8751 ( .ip1(n11060), .ip2(n10870), .op(n8638) );
  nand2_1 U8752 ( .ip1(n12235), .ip2(\cache_data[10][69] ), .op(n8620) );
  nand2_1 U8753 ( .ip1(n8905), .ip2(\cache_data[6][69] ), .op(n8619) );
  nand2_1 U8754 ( .ip1(n12152), .ip2(\cache_data[9][69] ), .op(n8618) );
  nand2_1 U8755 ( .ip1(n9681), .ip2(\cache_data[15][69] ), .op(n8617) );
  nand4_1 U8756 ( .ip1(n8620), .ip2(n8619), .ip3(n8618), .ip4(n8617), .op(
        n8636) );
  nand2_1 U8757 ( .ip1(n8911), .ip2(\cache_data[0][69] ), .op(n8624) );
  nand2_1 U8758 ( .ip1(n8900), .ip2(\cache_data[2][69] ), .op(n8623) );
  nand2_1 U8759 ( .ip1(n12240), .ip2(\cache_data[5][69] ), .op(n8622) );
  nand2_1 U8760 ( .ip1(n12234), .ip2(\cache_data[8][69] ), .op(n8621) );
  nand4_1 U8761 ( .ip1(n8624), .ip2(n8623), .ip3(n8622), .ip4(n8621), .op(
        n8635) );
  nand2_1 U8762 ( .ip1(n8899), .ip2(\cache_data[13][69] ), .op(n8628) );
  nand2_1 U8763 ( .ip1(n8906), .ip2(\cache_data[4][69] ), .op(n8627) );
  nand2_1 U8764 ( .ip1(n9669), .ip2(\cache_data[11][69] ), .op(n8626) );
  nand2_1 U8765 ( .ip1(n12207), .ip2(\cache_data[12][69] ), .op(n8625) );
  nand4_1 U8766 ( .ip1(n8628), .ip2(n8627), .ip3(n8626), .ip4(n8625), .op(
        n8634) );
  nand2_1 U8767 ( .ip1(n8894), .ip2(\cache_data[1][69] ), .op(n8632) );
  nand2_1 U8768 ( .ip1(n11971), .ip2(\cache_data[14][69] ), .op(n8631) );
  nand2_1 U8769 ( .ip1(n12219), .ip2(\cache_data[3][69] ), .op(n8630) );
  nand2_1 U8770 ( .ip1(n9670), .ip2(\cache_data[7][69] ), .op(n8629) );
  nand4_1 U8771 ( .ip1(n8632), .ip2(n8631), .ip3(n8630), .ip4(n8629), .op(
        n8633) );
  nor4_1 U8772 ( .ip1(n8636), .ip2(n8635), .ip3(n8634), .ip4(n8633), .op(
        n11059) );
  nor2_1 U8773 ( .ip1(n11059), .ip2(n10849), .op(n8637) );
  not_ab_or_c_or_d U8774 ( .ip1(n10894), .ip2(n11058), .ip3(n8638), .ip4(n8637), .op(n8660) );
  nand2_1 U8775 ( .ip1(n12226), .ip2(\cache_data[7][5] ), .op(n8642) );
  nand2_1 U8776 ( .ip1(n10975), .ip2(\cache_data[15][5] ), .op(n8641) );
  nand2_1 U8777 ( .ip1(n12220), .ip2(\cache_data[14][5] ), .op(n8640) );
  nand2_1 U8778 ( .ip1(n8906), .ip2(\cache_data[4][5] ), .op(n8639) );
  nand4_1 U8779 ( .ip1(n8642), .ip2(n8641), .ip3(n8640), .ip4(n8639), .op(
        n8658) );
  nand2_1 U8780 ( .ip1(n8900), .ip2(\cache_data[2][5] ), .op(n8646) );
  nand2_1 U8781 ( .ip1(n8894), .ip2(\cache_data[1][5] ), .op(n8645) );
  nand2_1 U8782 ( .ip1(n8905), .ip2(\cache_data[6][5] ), .op(n8644) );
  nand2_1 U8783 ( .ip1(n12121), .ip2(\cache_data[8][5] ), .op(n8643) );
  nand4_1 U8784 ( .ip1(n8646), .ip2(n8645), .ip3(n8644), .ip4(n8643), .op(
        n8657) );
  nand2_1 U8785 ( .ip1(n12207), .ip2(\cache_data[12][5] ), .op(n8650) );
  nand2_1 U8786 ( .ip1(n10964), .ip2(\cache_data[5][5] ), .op(n8649) );
  nand2_1 U8787 ( .ip1(n11317), .ip2(\cache_data[3][5] ), .op(n8648) );
  nand2_1 U8788 ( .ip1(n12096), .ip2(\cache_data[11][5] ), .op(n8647) );
  nand4_1 U8789 ( .ip1(n8650), .ip2(n8649), .ip3(n8648), .ip4(n8647), .op(
        n8656) );
  nand2_1 U8790 ( .ip1(n12126), .ip2(\cache_data[9][5] ), .op(n8654) );
  nand2_1 U8791 ( .ip1(n8899), .ip2(\cache_data[13][5] ), .op(n8653) );
  nand2_1 U8792 ( .ip1(n12235), .ip2(\cache_data[10][5] ), .op(n8652) );
  nand2_1 U8793 ( .ip1(n8911), .ip2(\cache_data[0][5] ), .op(n8651) );
  nand4_1 U8794 ( .ip1(n8654), .ip2(n8653), .ip3(n8652), .ip4(n8651), .op(
        n8655) );
  or4_1 U8795 ( .ip1(n8658), .ip2(n8657), .ip3(n8656), .ip4(n8655), .op(n11063) );
  nand2_1 U8796 ( .ip1(n10828), .ip2(n11063), .op(n8659) );
  nand3_1 U8797 ( .ip1(n8661), .ip2(n8660), .ip3(n8659), .op(n7443) );
  nand2_1 U8798 ( .ip1(data_wr_mem[6]), .ip2(n10873), .op(n8746) );
  nand2_1 U8799 ( .ip1(n12191), .ip2(\cache_data[8][6] ), .op(n8665) );
  nand2_1 U8800 ( .ip1(n8905), .ip2(\cache_data[6][6] ), .op(n8664) );
  nand2_1 U8801 ( .ip1(n8906), .ip2(\cache_data[4][6] ), .op(n8663) );
  nand2_1 U8802 ( .ip1(n8911), .ip2(\cache_data[0][6] ), .op(n8662) );
  nand4_1 U8803 ( .ip1(n8665), .ip2(n8664), .ip3(n8663), .ip4(n8662), .op(
        n8681) );
  nand2_1 U8804 ( .ip1(n12221), .ip2(\cache_data[15][6] ), .op(n8669) );
  nand2_1 U8805 ( .ip1(n12202), .ip2(\cache_data[7][6] ), .op(n8668) );
  nand2_1 U8806 ( .ip1(n11971), .ip2(\cache_data[14][6] ), .op(n8667) );
  nand2_1 U8807 ( .ip1(n12207), .ip2(\cache_data[12][6] ), .op(n8666) );
  nand4_1 U8808 ( .ip1(n8669), .ip2(n8668), .ip3(n8667), .ip4(n8666), .op(
        n8680) );
  nand2_1 U8809 ( .ip1(n12235), .ip2(\cache_data[10][6] ), .op(n8673) );
  nand2_1 U8810 ( .ip1(n12096), .ip2(\cache_data[11][6] ), .op(n8672) );
  nand2_1 U8811 ( .ip1(n8899), .ip2(\cache_data[13][6] ), .op(n8671) );
  nand2_1 U8812 ( .ip1(n12120), .ip2(\cache_data[1][6] ), .op(n8670) );
  nand4_1 U8813 ( .ip1(n8673), .ip2(n8672), .ip3(n8671), .ip4(n8670), .op(
        n8679) );
  nand2_1 U8814 ( .ip1(n8900), .ip2(\cache_data[2][6] ), .op(n8677) );
  nand2_1 U8815 ( .ip1(n12126), .ip2(\cache_data[9][6] ), .op(n8676) );
  nand2_1 U8816 ( .ip1(n12219), .ip2(\cache_data[3][6] ), .op(n8675) );
  nand2_1 U8817 ( .ip1(n12240), .ip2(\cache_data[5][6] ), .op(n8674) );
  nand4_1 U8818 ( .ip1(n8677), .ip2(n8676), .ip3(n8675), .ip4(n8674), .op(
        n8678) );
  or4_1 U8819 ( .ip1(n8681), .ip2(n8680), .ip3(n8679), .ip4(n8678), .op(n11067) );
  nand2_1 U8820 ( .ip1(n12235), .ip2(\cache_data[10][38] ), .op(n8685) );
  nand2_1 U8821 ( .ip1(n8905), .ip2(\cache_data[6][38] ), .op(n8684) );
  nand2_1 U8822 ( .ip1(n8911), .ip2(\cache_data[0][38] ), .op(n8683) );
  nand2_1 U8823 ( .ip1(n8900), .ip2(\cache_data[2][38] ), .op(n8682) );
  nand4_1 U8824 ( .ip1(n8685), .ip2(n8684), .ip3(n8683), .ip4(n8682), .op(
        n8701) );
  nand2_1 U8825 ( .ip1(n11971), .ip2(\cache_data[14][38] ), .op(n8689) );
  nand2_1 U8826 ( .ip1(n8906), .ip2(\cache_data[4][38] ), .op(n8688) );
  nand2_1 U8827 ( .ip1(n12096), .ip2(\cache_data[11][38] ), .op(n8687) );
  nand2_1 U8828 ( .ip1(n12207), .ip2(\cache_data[12][38] ), .op(n8686) );
  nand4_1 U8829 ( .ip1(n8689), .ip2(n8688), .ip3(n8687), .ip4(n8686), .op(
        n8700) );
  nand2_1 U8830 ( .ip1(n12126), .ip2(\cache_data[9][38] ), .op(n8693) );
  nand2_1 U8831 ( .ip1(n12221), .ip2(\cache_data[15][38] ), .op(n8692) );
  nand2_1 U8832 ( .ip1(n8899), .ip2(\cache_data[13][38] ), .op(n8691) );
  nand2_1 U8833 ( .ip1(n9675), .ip2(\cache_data[5][38] ), .op(n8690) );
  nand4_1 U8834 ( .ip1(n8693), .ip2(n8692), .ip3(n8691), .ip4(n8690), .op(
        n8699) );
  nand2_1 U8835 ( .ip1(n8894), .ip2(\cache_data[1][38] ), .op(n8697) );
  nand2_1 U8836 ( .ip1(n12202), .ip2(\cache_data[7][38] ), .op(n8696) );
  nand2_1 U8837 ( .ip1(n12219), .ip2(\cache_data[3][38] ), .op(n8695) );
  nand2_1 U8838 ( .ip1(n9668), .ip2(\cache_data[8][38] ), .op(n8694) );
  nand4_1 U8839 ( .ip1(n8697), .ip2(n8696), .ip3(n8695), .ip4(n8694), .op(
        n8698) );
  nor4_1 U8840 ( .ip1(n8701), .ip2(n8700), .ip3(n8699), .ip4(n8698), .op(
        n11069) );
  nor2_1 U8841 ( .ip1(n11069), .ip2(n10870), .op(n8723) );
  nand2_1 U8842 ( .ip1(n12126), .ip2(\cache_data[9][70] ), .op(n8705) );
  nand2_1 U8843 ( .ip1(n8906), .ip2(\cache_data[4][70] ), .op(n8704) );
  nand2_1 U8844 ( .ip1(n12220), .ip2(\cache_data[14][70] ), .op(n8703) );
  nand2_1 U8845 ( .ip1(n11317), .ip2(\cache_data[3][70] ), .op(n8702) );
  nand4_1 U8846 ( .ip1(n8705), .ip2(n8704), .ip3(n8703), .ip4(n8702), .op(
        n8721) );
  nand2_1 U8847 ( .ip1(n12202), .ip2(\cache_data[7][70] ), .op(n8709) );
  nand2_1 U8848 ( .ip1(n8905), .ip2(\cache_data[6][70] ), .op(n8708) );
  nand2_1 U8849 ( .ip1(n12240), .ip2(\cache_data[5][70] ), .op(n8707) );
  nand2_1 U8850 ( .ip1(n9681), .ip2(\cache_data[15][70] ), .op(n8706) );
  nand4_1 U8851 ( .ip1(n8709), .ip2(n8708), .ip3(n8707), .ip4(n8706), .op(
        n8720) );
  nand2_1 U8852 ( .ip1(n12191), .ip2(\cache_data[8][70] ), .op(n8713) );
  nand2_1 U8853 ( .ip1(n11927), .ip2(\cache_data[11][70] ), .op(n8712) );
  nand2_1 U8854 ( .ip1(n8900), .ip2(\cache_data[2][70] ), .op(n8711) );
  nand2_1 U8855 ( .ip1(n12227), .ip2(\cache_data[12][70] ), .op(n8710) );
  nand4_1 U8856 ( .ip1(n8713), .ip2(n8712), .ip3(n8711), .ip4(n8710), .op(
        n8719) );
  nand2_1 U8857 ( .ip1(n8894), .ip2(\cache_data[1][70] ), .op(n8717) );
  nand2_1 U8858 ( .ip1(n8899), .ip2(\cache_data[13][70] ), .op(n8716) );
  nand2_1 U8859 ( .ip1(n8911), .ip2(\cache_data[0][70] ), .op(n8715) );
  nand2_1 U8860 ( .ip1(n12235), .ip2(\cache_data[10][70] ), .op(n8714) );
  nand4_1 U8861 ( .ip1(n8717), .ip2(n8716), .ip3(n8715), .ip4(n8714), .op(
        n8718) );
  nor4_1 U8862 ( .ip1(n8721), .ip2(n8720), .ip3(n8719), .ip4(n8718), .op(
        n11068) );
  nor2_1 U8863 ( .ip1(n11068), .ip2(n10849), .op(n8722) );
  not_ab_or_c_or_d U8864 ( .ip1(n10828), .ip2(n11067), .ip3(n8723), .ip4(n8722), .op(n8745) );
  nand2_1 U8865 ( .ip1(n12126), .ip2(\cache_data[9][102] ), .op(n8727) );
  nand2_1 U8866 ( .ip1(n12096), .ip2(\cache_data[11][102] ), .op(n8726) );
  nand2_1 U8867 ( .ip1(n12240), .ip2(\cache_data[5][102] ), .op(n8725) );
  nand2_1 U8868 ( .ip1(n12219), .ip2(\cache_data[3][102] ), .op(n8724) );
  nand4_1 U8869 ( .ip1(n8727), .ip2(n8726), .ip3(n8725), .ip4(n8724), .op(
        n8743) );
  nand2_1 U8870 ( .ip1(n11971), .ip2(\cache_data[14][102] ), .op(n8731) );
  nand2_1 U8871 ( .ip1(n8899), .ip2(\cache_data[13][102] ), .op(n8730) );
  nand2_1 U8872 ( .ip1(n12235), .ip2(\cache_data[10][102] ), .op(n8729) );
  nand2_1 U8873 ( .ip1(n12221), .ip2(\cache_data[15][102] ), .op(n8728) );
  nand4_1 U8874 ( .ip1(n8731), .ip2(n8730), .ip3(n8729), .ip4(n8728), .op(
        n8742) );
  nand2_1 U8875 ( .ip1(n8905), .ip2(\cache_data[6][102] ), .op(n8735) );
  nand2_1 U8876 ( .ip1(n8911), .ip2(\cache_data[0][102] ), .op(n8734) );
  nand2_1 U8877 ( .ip1(n12202), .ip2(\cache_data[7][102] ), .op(n8733) );
  nand2_1 U8878 ( .ip1(n12207), .ip2(\cache_data[12][102] ), .op(n8732) );
  nand4_1 U8879 ( .ip1(n8735), .ip2(n8734), .ip3(n8733), .ip4(n8732), .op(
        n8741) );
  nand2_1 U8880 ( .ip1(n8894), .ip2(\cache_data[1][102] ), .op(n8739) );
  nand2_1 U8881 ( .ip1(n8906), .ip2(\cache_data[4][102] ), .op(n8738) );
  nand2_1 U8882 ( .ip1(n8900), .ip2(\cache_data[2][102] ), .op(n8737) );
  nand2_1 U8883 ( .ip1(n12191), .ip2(\cache_data[8][102] ), .op(n8736) );
  nand4_1 U8884 ( .ip1(n8739), .ip2(n8738), .ip3(n8737), .ip4(n8736), .op(
        n8740) );
  or4_1 U8885 ( .ip1(n8743), .ip2(n8742), .ip3(n8741), .ip4(n8740), .op(n11072) );
  nand2_1 U8886 ( .ip1(n10894), .ip2(n11072), .op(n8744) );
  nand3_1 U8887 ( .ip1(n8746), .ip2(n8745), .ip3(n8744), .op(n7442) );
  nand2_1 U8888 ( .ip1(n12219), .ip2(\cache_data[3][7] ), .op(n8750) );
  nand2_1 U8889 ( .ip1(n12121), .ip2(\cache_data[8][7] ), .op(n8749) );
  nand2_1 U8890 ( .ip1(n8899), .ip2(\cache_data[13][7] ), .op(n8748) );
  nand2_1 U8891 ( .ip1(n8905), .ip2(\cache_data[6][7] ), .op(n8747) );
  nand4_1 U8892 ( .ip1(n8750), .ip2(n8749), .ip3(n8748), .ip4(n8747), .op(
        n8766) );
  nand2_1 U8893 ( .ip1(n12221), .ip2(\cache_data[15][7] ), .op(n8754) );
  nand2_1 U8894 ( .ip1(n8894), .ip2(\cache_data[1][7] ), .op(n8753) );
  nand2_1 U8895 ( .ip1(n12126), .ip2(\cache_data[9][7] ), .op(n8752) );
  nand2_1 U8896 ( .ip1(n12096), .ip2(\cache_data[11][7] ), .op(n8751) );
  nand4_1 U8897 ( .ip1(n8754), .ip2(n8753), .ip3(n8752), .ip4(n8751), .op(
        n8765) );
  nand2_1 U8898 ( .ip1(n8911), .ip2(\cache_data[0][7] ), .op(n8758) );
  nand2_1 U8899 ( .ip1(n8900), .ip2(\cache_data[2][7] ), .op(n8757) );
  nand2_1 U8900 ( .ip1(n12207), .ip2(\cache_data[12][7] ), .op(n8756) );
  nand2_1 U8901 ( .ip1(n8906), .ip2(\cache_data[4][7] ), .op(n8755) );
  nand4_1 U8902 ( .ip1(n8758), .ip2(n8757), .ip3(n8756), .ip4(n8755), .op(
        n8764) );
  nand2_1 U8903 ( .ip1(n12226), .ip2(\cache_data[7][7] ), .op(n8762) );
  nand2_1 U8904 ( .ip1(n12235), .ip2(\cache_data[10][7] ), .op(n8761) );
  nand2_1 U8905 ( .ip1(n12240), .ip2(\cache_data[5][7] ), .op(n8760) );
  nand2_1 U8906 ( .ip1(n11971), .ip2(\cache_data[14][7] ), .op(n8759) );
  nand4_1 U8907 ( .ip1(n8762), .ip2(n8761), .ip3(n8760), .ip4(n8759), .op(
        n8763) );
  or4_1 U8908 ( .ip1(n8766), .ip2(n8765), .ip3(n8764), .ip4(n8763), .op(n11076) );
  nand2_1 U8909 ( .ip1(n10828), .ip2(n11076), .op(n8831) );
  nand2_1 U8910 ( .ip1(n12221), .ip2(\cache_data[15][71] ), .op(n8770) );
  nand2_1 U8911 ( .ip1(n8911), .ip2(\cache_data[0][71] ), .op(n8769) );
  nand2_1 U8912 ( .ip1(n8900), .ip2(\cache_data[2][71] ), .op(n8768) );
  nand2_1 U8913 ( .ip1(n12126), .ip2(\cache_data[9][71] ), .op(n8767) );
  nand4_1 U8914 ( .ip1(n8770), .ip2(n8769), .ip3(n8768), .ip4(n8767), .op(
        n8786) );
  nand2_1 U8915 ( .ip1(n11971), .ip2(\cache_data[14][71] ), .op(n8774) );
  nand2_1 U8916 ( .ip1(n8906), .ip2(\cache_data[4][71] ), .op(n8773) );
  nand2_1 U8917 ( .ip1(n8894), .ip2(\cache_data[1][71] ), .op(n8772) );
  nand2_1 U8918 ( .ip1(n12191), .ip2(\cache_data[8][71] ), .op(n8771) );
  nand4_1 U8919 ( .ip1(n8774), .ip2(n8773), .ip3(n8772), .ip4(n8771), .op(
        n8785) );
  nand2_1 U8920 ( .ip1(n12207), .ip2(\cache_data[12][71] ), .op(n8778) );
  nand2_1 U8921 ( .ip1(n11317), .ip2(\cache_data[3][71] ), .op(n8777) );
  nand2_1 U8922 ( .ip1(n8905), .ip2(\cache_data[6][71] ), .op(n8776) );
  nand2_1 U8923 ( .ip1(n12235), .ip2(\cache_data[10][71] ), .op(n8775) );
  nand4_1 U8924 ( .ip1(n8778), .ip2(n8777), .ip3(n8776), .ip4(n8775), .op(
        n8784) );
  nand2_1 U8925 ( .ip1(n12240), .ip2(\cache_data[5][71] ), .op(n8782) );
  nand2_1 U8926 ( .ip1(n9669), .ip2(\cache_data[11][71] ), .op(n8781) );
  nand2_1 U8927 ( .ip1(n12202), .ip2(\cache_data[7][71] ), .op(n8780) );
  nand2_1 U8928 ( .ip1(n8899), .ip2(\cache_data[13][71] ), .op(n8779) );
  nand4_1 U8929 ( .ip1(n8782), .ip2(n8781), .ip3(n8780), .ip4(n8779), .op(
        n8783) );
  nor4_1 U8930 ( .ip1(n8786), .ip2(n8785), .ip3(n8784), .ip4(n8783), .op(
        n11077) );
  nor2_1 U8931 ( .ip1(n11077), .ip2(n10849), .op(n8808) );
  nand2_1 U8932 ( .ip1(n8900), .ip2(\cache_data[2][39] ), .op(n8790) );
  nand2_1 U8933 ( .ip1(n12096), .ip2(\cache_data[11][39] ), .op(n8789) );
  nand2_1 U8934 ( .ip1(n8894), .ip2(\cache_data[1][39] ), .op(n8788) );
  nand2_1 U8935 ( .ip1(n8905), .ip2(\cache_data[6][39] ), .op(n8787) );
  nand4_1 U8936 ( .ip1(n8790), .ip2(n8789), .ip3(n8788), .ip4(n8787), .op(
        n8806) );
  nand2_1 U8937 ( .ip1(n11971), .ip2(\cache_data[14][39] ), .op(n8794) );
  nand2_1 U8938 ( .ip1(n12241), .ip2(\cache_data[9][39] ), .op(n8793) );
  nand2_1 U8939 ( .ip1(n9681), .ip2(\cache_data[15][39] ), .op(n8792) );
  nand2_1 U8940 ( .ip1(n8899), .ip2(\cache_data[13][39] ), .op(n8791) );
  nand4_1 U8941 ( .ip1(n8794), .ip2(n8793), .ip3(n8792), .ip4(n8791), .op(
        n8805) );
  nand2_1 U8942 ( .ip1(n12207), .ip2(\cache_data[12][39] ), .op(n8798) );
  nand2_1 U8943 ( .ip1(n9675), .ip2(\cache_data[5][39] ), .op(n8797) );
  nand2_1 U8944 ( .ip1(n12219), .ip2(\cache_data[3][39] ), .op(n8796) );
  nand2_1 U8945 ( .ip1(n8906), .ip2(\cache_data[4][39] ), .op(n8795) );
  nand4_1 U8946 ( .ip1(n8798), .ip2(n8797), .ip3(n8796), .ip4(n8795), .op(
        n8804) );
  nand2_1 U8947 ( .ip1(n12202), .ip2(\cache_data[7][39] ), .op(n8802) );
  nand2_1 U8948 ( .ip1(n12234), .ip2(\cache_data[8][39] ), .op(n8801) );
  nand2_1 U8949 ( .ip1(n8911), .ip2(\cache_data[0][39] ), .op(n8800) );
  nand2_1 U8950 ( .ip1(n12196), .ip2(\cache_data[10][39] ), .op(n8799) );
  nand4_1 U8951 ( .ip1(n8802), .ip2(n8801), .ip3(n8800), .ip4(n8799), .op(
        n8803) );
  nor4_1 U8952 ( .ip1(n8806), .ip2(n8805), .ip3(n8804), .ip4(n8803), .op(
        n11078) );
  nor2_1 U8953 ( .ip1(n11078), .ip2(n10870), .op(n8807) );
  not_ab_or_c_or_d U8954 ( .ip1(data_wr_mem[7]), .ip2(n10873), .ip3(n8808), 
        .ip4(n8807), .op(n8830) );
  nand2_1 U8955 ( .ip1(n12207), .ip2(\cache_data[12][103] ), .op(n8812) );
  nand2_1 U8956 ( .ip1(n8899), .ip2(\cache_data[13][103] ), .op(n8811) );
  nand2_1 U8957 ( .ip1(n12191), .ip2(\cache_data[8][103] ), .op(n8810) );
  nand2_1 U8958 ( .ip1(n8911), .ip2(\cache_data[0][103] ), .op(n8809) );
  nand4_1 U8959 ( .ip1(n8812), .ip2(n8811), .ip3(n8810), .ip4(n8809), .op(
        n8828) );
  nand2_1 U8960 ( .ip1(n8894), .ip2(\cache_data[1][103] ), .op(n8816) );
  nand2_1 U8961 ( .ip1(n12221), .ip2(\cache_data[15][103] ), .op(n8815) );
  nand2_1 U8962 ( .ip1(n12202), .ip2(\cache_data[7][103] ), .op(n8814) );
  nand2_1 U8963 ( .ip1(n8900), .ip2(\cache_data[2][103] ), .op(n8813) );
  nand4_1 U8964 ( .ip1(n8816), .ip2(n8815), .ip3(n8814), .ip4(n8813), .op(
        n8827) );
  nand2_1 U8965 ( .ip1(n8906), .ip2(\cache_data[4][103] ), .op(n8820) );
  nand2_1 U8966 ( .ip1(n11971), .ip2(\cache_data[14][103] ), .op(n8819) );
  nand2_1 U8967 ( .ip1(n12096), .ip2(\cache_data[11][103] ), .op(n8818) );
  nand2_1 U8968 ( .ip1(n12240), .ip2(\cache_data[5][103] ), .op(n8817) );
  nand4_1 U8969 ( .ip1(n8820), .ip2(n8819), .ip3(n8818), .ip4(n8817), .op(
        n8826) );
  nand2_1 U8970 ( .ip1(n8905), .ip2(\cache_data[6][103] ), .op(n8824) );
  nand2_1 U8971 ( .ip1(n12235), .ip2(\cache_data[10][103] ), .op(n8823) );
  nand2_1 U8972 ( .ip1(n12126), .ip2(\cache_data[9][103] ), .op(n8822) );
  nand2_1 U8973 ( .ip1(n12219), .ip2(\cache_data[3][103] ), .op(n8821) );
  nand4_1 U8974 ( .ip1(n8824), .ip2(n8823), .ip3(n8822), .ip4(n8821), .op(
        n8825) );
  or4_1 U8975 ( .ip1(n8828), .ip2(n8827), .ip3(n8826), .ip4(n8825), .op(n11081) );
  nand2_1 U8976 ( .ip1(n10894), .ip2(n11081), .op(n8829) );
  nand3_1 U8977 ( .ip1(n8831), .ip2(n8830), .ip3(n8829), .op(n7441) );
  nand2_1 U8978 ( .ip1(n8899), .ip2(\cache_data[13][8] ), .op(n8835) );
  nand2_1 U8979 ( .ip1(n12207), .ip2(\cache_data[12][8] ), .op(n8834) );
  nand2_1 U8980 ( .ip1(n8894), .ip2(\cache_data[1][8] ), .op(n8833) );
  nand2_1 U8981 ( .ip1(n8905), .ip2(\cache_data[6][8] ), .op(n8832) );
  nand4_1 U8982 ( .ip1(n8835), .ip2(n8834), .ip3(n8833), .ip4(n8832), .op(
        n8851) );
  nand2_1 U8983 ( .ip1(n12221), .ip2(\cache_data[15][8] ), .op(n8839) );
  nand2_1 U8984 ( .ip1(n12126), .ip2(\cache_data[9][8] ), .op(n8838) );
  nand2_1 U8985 ( .ip1(n12096), .ip2(\cache_data[11][8] ), .op(n8837) );
  nand2_1 U8986 ( .ip1(n12226), .ip2(\cache_data[7][8] ), .op(n8836) );
  nand4_1 U8987 ( .ip1(n8839), .ip2(n8838), .ip3(n8837), .ip4(n8836), .op(
        n8850) );
  nand2_1 U8988 ( .ip1(n12235), .ip2(\cache_data[10][8] ), .op(n8843) );
  nand2_1 U8989 ( .ip1(n12240), .ip2(\cache_data[5][8] ), .op(n8842) );
  nand2_1 U8990 ( .ip1(n11971), .ip2(\cache_data[14][8] ), .op(n8841) );
  nand2_1 U8991 ( .ip1(n12121), .ip2(\cache_data[8][8] ), .op(n8840) );
  nand4_1 U8992 ( .ip1(n8843), .ip2(n8842), .ip3(n8841), .ip4(n8840), .op(
        n8849) );
  nand2_1 U8993 ( .ip1(n12219), .ip2(\cache_data[3][8] ), .op(n8847) );
  nand2_1 U8994 ( .ip1(n8900), .ip2(\cache_data[2][8] ), .op(n8846) );
  nand2_1 U8995 ( .ip1(n8906), .ip2(\cache_data[4][8] ), .op(n8845) );
  nand2_1 U8996 ( .ip1(n8911), .ip2(\cache_data[0][8] ), .op(n8844) );
  nand4_1 U8997 ( .ip1(n8847), .ip2(n8846), .ip3(n8845), .ip4(n8844), .op(
        n8848) );
  or4_1 U8998 ( .ip1(n8851), .ip2(n8850), .ip3(n8849), .ip4(n8848), .op(n11085) );
  nand2_1 U8999 ( .ip1(n10828), .ip2(n11085), .op(n8922) );
  nand2_1 U9000 ( .ip1(n8906), .ip2(\cache_data[4][40] ), .op(n8855) );
  nand2_1 U9001 ( .ip1(n12240), .ip2(\cache_data[5][40] ), .op(n8854) );
  nand2_1 U9002 ( .ip1(n12191), .ip2(\cache_data[8][40] ), .op(n8853) );
  nand2_1 U9003 ( .ip1(n12207), .ip2(\cache_data[12][40] ), .op(n8852) );
  nand4_1 U9004 ( .ip1(n8855), .ip2(n8854), .ip3(n8853), .ip4(n8852), .op(
        n8871) );
  nand2_1 U9005 ( .ip1(n8894), .ip2(\cache_data[1][40] ), .op(n8859) );
  nand2_1 U9006 ( .ip1(n12226), .ip2(\cache_data[7][40] ), .op(n8858) );
  nand2_1 U9007 ( .ip1(n12235), .ip2(\cache_data[10][40] ), .op(n8857) );
  nand2_1 U9008 ( .ip1(n12221), .ip2(\cache_data[15][40] ), .op(n8856) );
  nand4_1 U9009 ( .ip1(n8859), .ip2(n8858), .ip3(n8857), .ip4(n8856), .op(
        n8870) );
  nand2_1 U9010 ( .ip1(n12096), .ip2(\cache_data[11][40] ), .op(n8863) );
  nand2_1 U9011 ( .ip1(n12219), .ip2(\cache_data[3][40] ), .op(n8862) );
  nand2_1 U9012 ( .ip1(n8905), .ip2(\cache_data[6][40] ), .op(n8861) );
  nand2_1 U9013 ( .ip1(n8900), .ip2(\cache_data[2][40] ), .op(n8860) );
  nand4_1 U9014 ( .ip1(n8863), .ip2(n8862), .ip3(n8861), .ip4(n8860), .op(
        n8869) );
  nand2_1 U9015 ( .ip1(n11971), .ip2(\cache_data[14][40] ), .op(n8867) );
  nand2_1 U9016 ( .ip1(n12126), .ip2(\cache_data[9][40] ), .op(n8866) );
  nand2_1 U9017 ( .ip1(n8911), .ip2(\cache_data[0][40] ), .op(n8865) );
  nand2_1 U9018 ( .ip1(n8899), .ip2(\cache_data[13][40] ), .op(n8864) );
  nand4_1 U9019 ( .ip1(n8867), .ip2(n8866), .ip3(n8865), .ip4(n8864), .op(
        n8868) );
  nor4_1 U9020 ( .ip1(n8871), .ip2(n8870), .ip3(n8869), .ip4(n8868), .op(
        n11087) );
  nor2_1 U9021 ( .ip1(n11087), .ip2(n10870), .op(n8893) );
  nand2_1 U9022 ( .ip1(n8905), .ip2(\cache_data[6][72] ), .op(n8875) );
  nand2_1 U9023 ( .ip1(n8911), .ip2(\cache_data[0][72] ), .op(n8874) );
  nand2_1 U9024 ( .ip1(n8899), .ip2(\cache_data[13][72] ), .op(n8873) );
  nand2_1 U9025 ( .ip1(n12120), .ip2(\cache_data[1][72] ), .op(n8872) );
  nand4_1 U9026 ( .ip1(n8875), .ip2(n8874), .ip3(n8873), .ip4(n8872), .op(
        n8891) );
  nand2_1 U9027 ( .ip1(n12096), .ip2(\cache_data[11][72] ), .op(n8879) );
  nand2_1 U9028 ( .ip1(n12202), .ip2(\cache_data[7][72] ), .op(n8878) );
  nand2_1 U9029 ( .ip1(n12191), .ip2(\cache_data[8][72] ), .op(n8877) );
  nand2_1 U9030 ( .ip1(n12207), .ip2(\cache_data[12][72] ), .op(n8876) );
  nand4_1 U9031 ( .ip1(n8879), .ip2(n8878), .ip3(n8877), .ip4(n8876), .op(
        n8890) );
  nand2_1 U9032 ( .ip1(n12219), .ip2(\cache_data[3][72] ), .op(n8883) );
  nand2_1 U9033 ( .ip1(n12126), .ip2(\cache_data[9][72] ), .op(n8882) );
  nand2_1 U9034 ( .ip1(n12221), .ip2(\cache_data[15][72] ), .op(n8881) );
  nand2_1 U9035 ( .ip1(n12240), .ip2(\cache_data[5][72] ), .op(n8880) );
  nand4_1 U9036 ( .ip1(n8883), .ip2(n8882), .ip3(n8881), .ip4(n8880), .op(
        n8889) );
  nand2_1 U9037 ( .ip1(n8906), .ip2(\cache_data[4][72] ), .op(n8887) );
  nand2_1 U9038 ( .ip1(n12220), .ip2(\cache_data[14][72] ), .op(n8886) );
  nand2_1 U9039 ( .ip1(n8900), .ip2(\cache_data[2][72] ), .op(n8885) );
  nand2_1 U9040 ( .ip1(n12235), .ip2(\cache_data[10][72] ), .op(n8884) );
  nand4_1 U9041 ( .ip1(n8887), .ip2(n8886), .ip3(n8885), .ip4(n8884), .op(
        n8888) );
  nor4_1 U9042 ( .ip1(n8891), .ip2(n8890), .ip3(n8889), .ip4(n8888), .op(
        n11086) );
  nor2_1 U9043 ( .ip1(n11086), .ip2(n10849), .op(n8892) );
  not_ab_or_c_or_d U9044 ( .ip1(data_wr_mem[8]), .ip2(n10873), .ip3(n8893), 
        .ip4(n8892), .op(n8921) );
  nand2_1 U9045 ( .ip1(n8894), .ip2(\cache_data[1][104] ), .op(n8898) );
  nand2_1 U9046 ( .ip1(n12126), .ip2(\cache_data[9][104] ), .op(n8897) );
  nand2_1 U9047 ( .ip1(n12221), .ip2(\cache_data[15][104] ), .op(n8896) );
  nand2_1 U9048 ( .ip1(n12219), .ip2(\cache_data[3][104] ), .op(n8895) );
  nand4_1 U9049 ( .ip1(n8898), .ip2(n8897), .ip3(n8896), .ip4(n8895), .op(
        n8919) );
  nand2_1 U9050 ( .ip1(n8899), .ip2(\cache_data[13][104] ), .op(n8904) );
  nand2_1 U9051 ( .ip1(n12096), .ip2(\cache_data[11][104] ), .op(n8903) );
  nand2_1 U9052 ( .ip1(n8900), .ip2(\cache_data[2][104] ), .op(n8902) );
  nand2_1 U9053 ( .ip1(n12240), .ip2(\cache_data[5][104] ), .op(n8901) );
  nand4_1 U9054 ( .ip1(n8904), .ip2(n8903), .ip3(n8902), .ip4(n8901), .op(
        n8918) );
  nand2_1 U9055 ( .ip1(n8905), .ip2(\cache_data[6][104] ), .op(n8910) );
  nand2_1 U9056 ( .ip1(n12235), .ip2(\cache_data[10][104] ), .op(n8909) );
  nand2_1 U9057 ( .ip1(n8906), .ip2(\cache_data[4][104] ), .op(n8908) );
  nand2_1 U9058 ( .ip1(n12207), .ip2(\cache_data[12][104] ), .op(n8907) );
  nand4_1 U9059 ( .ip1(n8910), .ip2(n8909), .ip3(n8908), .ip4(n8907), .op(
        n8917) );
  nand2_1 U9060 ( .ip1(n11971), .ip2(\cache_data[14][104] ), .op(n8915) );
  nand2_1 U9061 ( .ip1(n12226), .ip2(\cache_data[7][104] ), .op(n8914) );
  nand2_1 U9062 ( .ip1(n8911), .ip2(\cache_data[0][104] ), .op(n8913) );
  nand2_1 U9063 ( .ip1(n12121), .ip2(\cache_data[8][104] ), .op(n8912) );
  nand4_1 U9064 ( .ip1(n8915), .ip2(n8914), .ip3(n8913), .ip4(n8912), .op(
        n8916) );
  or4_1 U9065 ( .ip1(n8919), .ip2(n8918), .ip3(n8917), .ip4(n8916), .op(n11090) );
  nand2_1 U9066 ( .ip1(n10894), .ip2(n11090), .op(n8920) );
  nand3_1 U9067 ( .ip1(n8922), .ip2(n8921), .ip3(n8920), .op(n7440) );
  nand2_1 U9068 ( .ip1(data_wr_mem[9]), .ip2(n10873), .op(n9009) );
  nand2_1 U9069 ( .ip1(n12201), .ip2(\cache_data[4][105] ), .op(n8927) );
  inv_1 U9070 ( .ip(n12233), .op(n8923) );
  inv_1 U9071 ( .ip(n8923), .op(n9688) );
  nand2_1 U9072 ( .ip1(n9688), .ip2(\cache_data[0][105] ), .op(n8926) );
  inv_1 U9073 ( .ip(n11612), .op(n9681) );
  nand2_1 U9074 ( .ip1(n9681), .ip2(\cache_data[15][105] ), .op(n8925) );
  nand2_1 U9075 ( .ip1(n12179), .ip2(\cache_data[6][105] ), .op(n8924) );
  nand4_1 U9076 ( .ip1(n8927), .ip2(n8926), .ip3(n8925), .ip4(n8924), .op(
        n8944) );
  inv_1 U9077 ( .ip(n8144), .op(n9682) );
  nand2_1 U9078 ( .ip1(n9682), .ip2(\cache_data[9][105] ), .op(n8932) );
  nand2_1 U9079 ( .ip1(n12165), .ip2(\cache_data[13][105] ), .op(n8931) );
  inv_1 U9080 ( .ip(n8137), .op(n9668) );
  nand2_1 U9081 ( .ip1(n9668), .ip2(\cache_data[8][105] ), .op(n8930) );
  inv_1 U9082 ( .ip(n12228), .op(n8928) );
  inv_1 U9083 ( .ip(n8928), .op(n9687) );
  nand2_1 U9084 ( .ip1(n9687), .ip2(\cache_data[2][105] ), .op(n8929) );
  nand4_1 U9085 ( .ip1(n8932), .ip2(n8931), .ip3(n8930), .ip4(n8929), .op(
        n8943) );
  inv_1 U9086 ( .ip(n11476), .op(n9680) );
  nand2_1 U9087 ( .ip1(n9680), .ip2(\cache_data[3][105] ), .op(n8936) );
  inv_1 U9088 ( .ip(n11600), .op(n9690) );
  nand2_1 U9089 ( .ip1(n9690), .ip2(\cache_data[14][105] ), .op(n8935) );
  nand2_1 U9090 ( .ip1(n11927), .ip2(\cache_data[11][105] ), .op(n8934) );
  inv_1 U9091 ( .ip(n11493), .op(n9675) );
  nand2_1 U9092 ( .ip1(n9675), .ip2(\cache_data[5][105] ), .op(n8933) );
  nand4_1 U9093 ( .ip1(n8936), .ip2(n8935), .ip3(n8934), .ip4(n8933), .op(
        n8942) );
  inv_1 U9094 ( .ip(n8146), .op(n9689) );
  nand2_1 U9095 ( .ip1(n9689), .ip2(\cache_data[10][105] ), .op(n8940) );
  nand2_1 U9096 ( .ip1(n12120), .ip2(\cache_data[1][105] ), .op(n8939) );
  inv_1 U9097 ( .ip(n8153), .op(n9670) );
  nand2_1 U9098 ( .ip1(n9670), .ip2(\cache_data[7][105] ), .op(n8938) );
  inv_1 U9099 ( .ip(n11551), .op(n9560) );
  nand2_1 U9100 ( .ip1(n9560), .ip2(\cache_data[12][105] ), .op(n8937) );
  nand4_1 U9101 ( .ip1(n8940), .ip2(n8939), .ip3(n8938), .ip4(n8937), .op(
        n8941) );
  or4_1 U9102 ( .ip1(n8944), .ip2(n8943), .ip3(n8942), .ip4(n8941), .op(n11094) );
  nand2_1 U9103 ( .ip1(n9668), .ip2(\cache_data[8][73] ), .op(n8948) );
  nand2_1 U9104 ( .ip1(n9689), .ip2(\cache_data[10][73] ), .op(n8947) );
  nand2_1 U9105 ( .ip1(n9682), .ip2(\cache_data[9][73] ), .op(n8946) );
  nand2_1 U9106 ( .ip1(n9560), .ip2(\cache_data[12][73] ), .op(n8945) );
  nand4_1 U9107 ( .ip1(n8948), .ip2(n8947), .ip3(n8946), .ip4(n8945), .op(
        n8964) );
  nand2_1 U9108 ( .ip1(n9690), .ip2(\cache_data[14][73] ), .op(n8952) );
  nand2_1 U9109 ( .ip1(n9688), .ip2(\cache_data[0][73] ), .op(n8951) );
  nand2_1 U9110 ( .ip1(n9670), .ip2(\cache_data[7][73] ), .op(n8950) );
  nand2_1 U9111 ( .ip1(n9681), .ip2(\cache_data[15][73] ), .op(n8949) );
  nand4_1 U9112 ( .ip1(n8952), .ip2(n8951), .ip3(n8950), .ip4(n8949), .op(
        n8963) );
  nand2_1 U9113 ( .ip1(n8905), .ip2(\cache_data[6][73] ), .op(n8956) );
  nand2_1 U9114 ( .ip1(n11927), .ip2(\cache_data[11][73] ), .op(n8955) );
  nand2_1 U9115 ( .ip1(n9687), .ip2(\cache_data[2][73] ), .op(n8954) );
  nand2_1 U9116 ( .ip1(n12120), .ip2(\cache_data[1][73] ), .op(n8953) );
  nand4_1 U9117 ( .ip1(n8956), .ip2(n8955), .ip3(n8954), .ip4(n8953), .op(
        n8962) );
  nand2_1 U9118 ( .ip1(n12142), .ip2(\cache_data[13][73] ), .op(n8960) );
  nand2_1 U9119 ( .ip1(n12164), .ip2(\cache_data[4][73] ), .op(n8959) );
  nand2_1 U9120 ( .ip1(n9680), .ip2(\cache_data[3][73] ), .op(n8958) );
  nand2_1 U9121 ( .ip1(n9675), .ip2(\cache_data[5][73] ), .op(n8957) );
  nand4_1 U9122 ( .ip1(n8960), .ip2(n8959), .ip3(n8958), .ip4(n8957), .op(
        n8961) );
  nor4_1 U9123 ( .ip1(n8964), .ip2(n8963), .ip3(n8962), .ip4(n8961), .op(
        n11095) );
  nor2_1 U9124 ( .ip1(n11095), .ip2(n10849), .op(n8986) );
  nand2_1 U9125 ( .ip1(n9682), .ip2(\cache_data[9][41] ), .op(n8968) );
  nand2_1 U9126 ( .ip1(n9668), .ip2(\cache_data[8][41] ), .op(n8967) );
  nand2_1 U9127 ( .ip1(n12120), .ip2(\cache_data[1][41] ), .op(n8966) );
  nand2_1 U9128 ( .ip1(n9688), .ip2(\cache_data[0][41] ), .op(n8965) );
  nand4_1 U9129 ( .ip1(n8968), .ip2(n8967), .ip3(n8966), .ip4(n8965), .op(
        n8984) );
  nand2_1 U9130 ( .ip1(n9690), .ip2(\cache_data[14][41] ), .op(n8972) );
  nand2_1 U9131 ( .ip1(n11927), .ip2(\cache_data[11][41] ), .op(n8971) );
  nand2_1 U9132 ( .ip1(n9681), .ip2(\cache_data[15][41] ), .op(n8970) );
  nand2_1 U9133 ( .ip1(n9687), .ip2(\cache_data[2][41] ), .op(n8969) );
  nand4_1 U9134 ( .ip1(n8972), .ip2(n8971), .ip3(n8970), .ip4(n8969), .op(
        n8983) );
  nand2_1 U9135 ( .ip1(n9675), .ip2(\cache_data[5][41] ), .op(n8976) );
  nand2_1 U9136 ( .ip1(n9670), .ip2(\cache_data[7][41] ), .op(n8975) );
  nand2_1 U9137 ( .ip1(n9560), .ip2(\cache_data[12][41] ), .op(n8974) );
  nand2_1 U9138 ( .ip1(n9689), .ip2(\cache_data[10][41] ), .op(n8973) );
  nand4_1 U9139 ( .ip1(n8976), .ip2(n8975), .ip3(n8974), .ip4(n8973), .op(
        n8982) );
  nand2_1 U9140 ( .ip1(n8905), .ip2(\cache_data[6][41] ), .op(n8980) );
  nand2_1 U9141 ( .ip1(n9680), .ip2(\cache_data[3][41] ), .op(n8979) );
  nand2_1 U9142 ( .ip1(n8899), .ip2(\cache_data[13][41] ), .op(n8978) );
  nand2_1 U9143 ( .ip1(n12243), .ip2(\cache_data[4][41] ), .op(n8977) );
  nand4_1 U9144 ( .ip1(n8980), .ip2(n8979), .ip3(n8978), .ip4(n8977), .op(
        n8981) );
  nor4_1 U9145 ( .ip1(n8984), .ip2(n8983), .ip3(n8982), .ip4(n8981), .op(
        n11096) );
  nor2_1 U9146 ( .ip1(n11096), .ip2(n10870), .op(n8985) );
  not_ab_or_c_or_d U9147 ( .ip1(n10894), .ip2(n11094), .ip3(n8986), .ip4(n8985), .op(n9008) );
  nand2_1 U9148 ( .ip1(n9682), .ip2(\cache_data[9][9] ), .op(n8990) );
  nand2_1 U9149 ( .ip1(n11927), .ip2(\cache_data[11][9] ), .op(n8989) );
  nand2_1 U9150 ( .ip1(n9675), .ip2(\cache_data[5][9] ), .op(n8988) );
  nand2_1 U9151 ( .ip1(n9687), .ip2(\cache_data[2][9] ), .op(n8987) );
  nand4_1 U9152 ( .ip1(n8990), .ip2(n8989), .ip3(n8988), .ip4(n8987), .op(
        n9006) );
  nand2_1 U9153 ( .ip1(n9680), .ip2(\cache_data[3][9] ), .op(n8994) );
  nand2_1 U9154 ( .ip1(n12165), .ip2(\cache_data[13][9] ), .op(n8993) );
  nand2_1 U9155 ( .ip1(n9681), .ip2(\cache_data[15][9] ), .op(n8992) );
  nand2_1 U9156 ( .ip1(n9690), .ip2(\cache_data[14][9] ), .op(n8991) );
  nand4_1 U9157 ( .ip1(n8994), .ip2(n8993), .ip3(n8992), .ip4(n8991), .op(
        n9005) );
  nand2_1 U9158 ( .ip1(n12201), .ip2(\cache_data[4][9] ), .op(n8998) );
  nand2_1 U9159 ( .ip1(n9689), .ip2(\cache_data[10][9] ), .op(n8997) );
  nand2_1 U9160 ( .ip1(n9668), .ip2(\cache_data[8][9] ), .op(n8996) );
  nand2_1 U9161 ( .ip1(n12120), .ip2(\cache_data[1][9] ), .op(n8995) );
  nand4_1 U9162 ( .ip1(n8998), .ip2(n8997), .ip3(n8996), .ip4(n8995), .op(
        n9004) );
  nand2_1 U9163 ( .ip1(n9688), .ip2(\cache_data[0][9] ), .op(n9002) );
  nand2_1 U9164 ( .ip1(n12179), .ip2(\cache_data[6][9] ), .op(n9001) );
  nand2_1 U9165 ( .ip1(n9670), .ip2(\cache_data[7][9] ), .op(n9000) );
  nand2_1 U9166 ( .ip1(n9560), .ip2(\cache_data[12][9] ), .op(n8999) );
  nand4_1 U9167 ( .ip1(n9002), .ip2(n9001), .ip3(n9000), .ip4(n8999), .op(
        n9003) );
  or4_1 U9168 ( .ip1(n9006), .ip2(n9005), .ip3(n9004), .ip4(n9003), .op(n11099) );
  nand2_1 U9169 ( .ip1(n10828), .ip2(n11099), .op(n9007) );
  nand3_1 U9170 ( .ip1(n9009), .ip2(n9008), .ip3(n9007), .op(n7439) );
  nand2_1 U9171 ( .ip1(n9682), .ip2(\cache_data[9][10] ), .op(n9013) );
  nand2_1 U9172 ( .ip1(n9668), .ip2(\cache_data[8][10] ), .op(n9012) );
  nand2_1 U9173 ( .ip1(n12096), .ip2(\cache_data[11][10] ), .op(n9011) );
  nand2_1 U9174 ( .ip1(n9690), .ip2(\cache_data[14][10] ), .op(n9010) );
  nand4_1 U9175 ( .ip1(n9013), .ip2(n9012), .ip3(n9011), .ip4(n9010), .op(
        n9029) );
  nand2_1 U9176 ( .ip1(n12120), .ip2(\cache_data[1][10] ), .op(n9017) );
  nand2_1 U9177 ( .ip1(n12142), .ip2(\cache_data[13][10] ), .op(n9016) );
  nand2_1 U9178 ( .ip1(n9687), .ip2(\cache_data[2][10] ), .op(n9015) );
  nand2_1 U9179 ( .ip1(n9560), .ip2(\cache_data[12][10] ), .op(n9014) );
  nand4_1 U9180 ( .ip1(n9017), .ip2(n9016), .ip3(n9015), .ip4(n9014), .op(
        n9028) );
  nand2_1 U9181 ( .ip1(n9689), .ip2(\cache_data[10][10] ), .op(n9021) );
  nand2_1 U9182 ( .ip1(n10305), .ip2(\cache_data[6][10] ), .op(n9020) );
  nand2_1 U9183 ( .ip1(n9688), .ip2(\cache_data[0][10] ), .op(n9019) );
  nand2_1 U9184 ( .ip1(n9681), .ip2(\cache_data[15][10] ), .op(n9018) );
  nand4_1 U9185 ( .ip1(n9021), .ip2(n9020), .ip3(n9019), .ip4(n9018), .op(
        n9027) );
  nand2_1 U9186 ( .ip1(n9675), .ip2(\cache_data[5][10] ), .op(n9025) );
  nand2_1 U9187 ( .ip1(n12201), .ip2(\cache_data[4][10] ), .op(n9024) );
  nand2_1 U9188 ( .ip1(n9670), .ip2(\cache_data[7][10] ), .op(n9023) );
  nand2_1 U9189 ( .ip1(n9680), .ip2(\cache_data[3][10] ), .op(n9022) );
  nand4_1 U9190 ( .ip1(n9025), .ip2(n9024), .ip3(n9023), .ip4(n9022), .op(
        n9026) );
  or4_1 U9191 ( .ip1(n9029), .ip2(n9028), .ip3(n9027), .ip4(n9026), .op(n11103) );
  nand2_1 U9192 ( .ip1(n10828), .ip2(n11103), .op(n9094) );
  nand2_1 U9193 ( .ip1(n12165), .ip2(\cache_data[13][42] ), .op(n9033) );
  nand2_1 U9194 ( .ip1(n9675), .ip2(\cache_data[5][42] ), .op(n9032) );
  nand2_1 U9195 ( .ip1(n11927), .ip2(\cache_data[11][42] ), .op(n9031) );
  nand2_1 U9196 ( .ip1(n12120), .ip2(\cache_data[1][42] ), .op(n9030) );
  nand4_1 U9197 ( .ip1(n9033), .ip2(n9032), .ip3(n9031), .ip4(n9030), .op(
        n9049) );
  nand2_1 U9198 ( .ip1(n9681), .ip2(\cache_data[15][42] ), .op(n9037) );
  nand2_1 U9199 ( .ip1(n9688), .ip2(\cache_data[0][42] ), .op(n9036) );
  nand2_1 U9200 ( .ip1(n9680), .ip2(\cache_data[3][42] ), .op(n9035) );
  nand2_1 U9201 ( .ip1(n9690), .ip2(\cache_data[14][42] ), .op(n9034) );
  nand4_1 U9202 ( .ip1(n9037), .ip2(n9036), .ip3(n9035), .ip4(n9034), .op(
        n9048) );
  nand2_1 U9203 ( .ip1(n9689), .ip2(\cache_data[10][42] ), .op(n9041) );
  nand2_1 U9204 ( .ip1(n12201), .ip2(\cache_data[4][42] ), .op(n9040) );
  nand2_1 U9205 ( .ip1(n9668), .ip2(\cache_data[8][42] ), .op(n9039) );
  nand2_1 U9206 ( .ip1(n9670), .ip2(\cache_data[7][42] ), .op(n9038) );
  nand4_1 U9207 ( .ip1(n9041), .ip2(n9040), .ip3(n9039), .ip4(n9038), .op(
        n9047) );
  nand2_1 U9208 ( .ip1(n9682), .ip2(\cache_data[9][42] ), .op(n9045) );
  nand2_1 U9209 ( .ip1(n10305), .ip2(\cache_data[6][42] ), .op(n9044) );
  nand2_1 U9210 ( .ip1(n9687), .ip2(\cache_data[2][42] ), .op(n9043) );
  nand2_1 U9211 ( .ip1(n9560), .ip2(\cache_data[12][42] ), .op(n9042) );
  nand4_1 U9212 ( .ip1(n9045), .ip2(n9044), .ip3(n9043), .ip4(n9042), .op(
        n9046) );
  nor4_1 U9213 ( .ip1(n9049), .ip2(n9048), .ip3(n9047), .ip4(n9046), .op(
        n11105) );
  nor2_1 U9214 ( .ip1(n11105), .ip2(n10870), .op(n9071) );
  nand2_1 U9215 ( .ip1(n12201), .ip2(\cache_data[4][74] ), .op(n9053) );
  nand2_1 U9216 ( .ip1(n12165), .ip2(\cache_data[13][74] ), .op(n9052) );
  nand2_1 U9217 ( .ip1(n9670), .ip2(\cache_data[7][74] ), .op(n9051) );
  nand2_1 U9218 ( .ip1(n8905), .ip2(\cache_data[6][74] ), .op(n9050) );
  nand4_1 U9219 ( .ip1(n9053), .ip2(n9052), .ip3(n9051), .ip4(n9050), .op(
        n9069) );
  nand2_1 U9220 ( .ip1(n9690), .ip2(\cache_data[14][74] ), .op(n9057) );
  nand2_1 U9221 ( .ip1(n12120), .ip2(\cache_data[1][74] ), .op(n9056) );
  nand2_1 U9222 ( .ip1(n9680), .ip2(\cache_data[3][74] ), .op(n9055) );
  nand2_1 U9223 ( .ip1(n11927), .ip2(\cache_data[11][74] ), .op(n9054) );
  nand4_1 U9224 ( .ip1(n9057), .ip2(n9056), .ip3(n9055), .ip4(n9054), .op(
        n9068) );
  nand2_1 U9225 ( .ip1(n9687), .ip2(\cache_data[2][74] ), .op(n9061) );
  nand2_1 U9226 ( .ip1(n9681), .ip2(\cache_data[15][74] ), .op(n9060) );
  nand2_1 U9227 ( .ip1(n9668), .ip2(\cache_data[8][74] ), .op(n9059) );
  nand2_1 U9228 ( .ip1(n9675), .ip2(\cache_data[5][74] ), .op(n9058) );
  nand4_1 U9229 ( .ip1(n9061), .ip2(n9060), .ip3(n9059), .ip4(n9058), .op(
        n9067) );
  nand2_1 U9230 ( .ip1(n9689), .ip2(\cache_data[10][74] ), .op(n9065) );
  nand2_1 U9231 ( .ip1(n9688), .ip2(\cache_data[0][74] ), .op(n9064) );
  nand2_1 U9232 ( .ip1(n9682), .ip2(\cache_data[9][74] ), .op(n9063) );
  nand2_1 U9233 ( .ip1(n9560), .ip2(\cache_data[12][74] ), .op(n9062) );
  nand4_1 U9234 ( .ip1(n9065), .ip2(n9064), .ip3(n9063), .ip4(n9062), .op(
        n9066) );
  nor4_1 U9235 ( .ip1(n9069), .ip2(n9068), .ip3(n9067), .ip4(n9066), .op(
        n11104) );
  nor2_1 U9236 ( .ip1(n11104), .ip2(n10849), .op(n9070) );
  not_ab_or_c_or_d U9237 ( .ip1(data_wr_mem[10]), .ip2(n10873), .ip3(n9071), 
        .ip4(n9070), .op(n9093) );
  nand2_1 U9238 ( .ip1(n9687), .ip2(\cache_data[2][106] ), .op(n9075) );
  nand2_1 U9239 ( .ip1(n9689), .ip2(\cache_data[10][106] ), .op(n9074) );
  nand2_1 U9240 ( .ip1(n9675), .ip2(\cache_data[5][106] ), .op(n9073) );
  nand2_1 U9241 ( .ip1(n12120), .ip2(\cache_data[1][106] ), .op(n9072) );
  nand4_1 U9242 ( .ip1(n9075), .ip2(n9074), .ip3(n9073), .ip4(n9072), .op(
        n9091) );
  nand2_1 U9243 ( .ip1(n9560), .ip2(\cache_data[12][106] ), .op(n9079) );
  nand2_1 U9244 ( .ip1(n9668), .ip2(\cache_data[8][106] ), .op(n9078) );
  nand2_1 U9245 ( .ip1(n12142), .ip2(\cache_data[13][106] ), .op(n9077) );
  nand2_1 U9246 ( .ip1(n10305), .ip2(\cache_data[6][106] ), .op(n9076) );
  nand4_1 U9247 ( .ip1(n9079), .ip2(n9078), .ip3(n9077), .ip4(n9076), .op(
        n9090) );
  nand2_1 U9248 ( .ip1(n12201), .ip2(\cache_data[4][106] ), .op(n9083) );
  nand2_1 U9249 ( .ip1(n9682), .ip2(\cache_data[9][106] ), .op(n9082) );
  nand2_1 U9250 ( .ip1(n12096), .ip2(\cache_data[11][106] ), .op(n9081) );
  nand2_1 U9251 ( .ip1(n9681), .ip2(\cache_data[15][106] ), .op(n9080) );
  nand4_1 U9252 ( .ip1(n9083), .ip2(n9082), .ip3(n9081), .ip4(n9080), .op(
        n9089) );
  nand2_1 U9253 ( .ip1(n9680), .ip2(\cache_data[3][106] ), .op(n9087) );
  nand2_1 U9254 ( .ip1(n9688), .ip2(\cache_data[0][106] ), .op(n9086) );
  nand2_1 U9255 ( .ip1(n9670), .ip2(\cache_data[7][106] ), .op(n9085) );
  nand2_1 U9256 ( .ip1(n9690), .ip2(\cache_data[14][106] ), .op(n9084) );
  nand4_1 U9257 ( .ip1(n9087), .ip2(n9086), .ip3(n9085), .ip4(n9084), .op(
        n9088) );
  or4_1 U9258 ( .ip1(n9091), .ip2(n9090), .ip3(n9089), .ip4(n9088), .op(n11108) );
  nand2_1 U9259 ( .ip1(n10894), .ip2(n11108), .op(n9092) );
  nand3_1 U9260 ( .ip1(n9094), .ip2(n9093), .ip3(n9092), .op(n7438) );
  nand2_1 U9261 ( .ip1(n12142), .ip2(\cache_data[13][11] ), .op(n9098) );
  nand2_1 U9262 ( .ip1(n9682), .ip2(\cache_data[9][11] ), .op(n9097) );
  nand2_1 U9263 ( .ip1(n9680), .ip2(\cache_data[3][11] ), .op(n9096) );
  nand2_1 U9264 ( .ip1(n9675), .ip2(\cache_data[5][11] ), .op(n9095) );
  nand4_1 U9265 ( .ip1(n9098), .ip2(n9097), .ip3(n9096), .ip4(n9095), .op(
        n9114) );
  nand2_1 U9266 ( .ip1(n9670), .ip2(\cache_data[7][11] ), .op(n9102) );
  nand2_1 U9267 ( .ip1(n9687), .ip2(\cache_data[2][11] ), .op(n9101) );
  nand2_1 U9268 ( .ip1(n12096), .ip2(\cache_data[11][11] ), .op(n9100) );
  nand2_1 U9269 ( .ip1(n9560), .ip2(\cache_data[12][11] ), .op(n9099) );
  nand4_1 U9270 ( .ip1(n9102), .ip2(n9101), .ip3(n9100), .ip4(n9099), .op(
        n9113) );
  nand2_1 U9271 ( .ip1(n9689), .ip2(\cache_data[10][11] ), .op(n9106) );
  nand2_1 U9272 ( .ip1(n9690), .ip2(\cache_data[14][11] ), .op(n9105) );
  nand2_1 U9273 ( .ip1(n12201), .ip2(\cache_data[4][11] ), .op(n9104) );
  nand2_1 U9274 ( .ip1(n10305), .ip2(\cache_data[6][11] ), .op(n9103) );
  nand4_1 U9275 ( .ip1(n9106), .ip2(n9105), .ip3(n9104), .ip4(n9103), .op(
        n9112) );
  nand2_1 U9276 ( .ip1(n9688), .ip2(\cache_data[0][11] ), .op(n9110) );
  nand2_1 U9277 ( .ip1(n9668), .ip2(\cache_data[8][11] ), .op(n9109) );
  nand2_1 U9278 ( .ip1(n9681), .ip2(\cache_data[15][11] ), .op(n9108) );
  nand2_1 U9279 ( .ip1(n12120), .ip2(\cache_data[1][11] ), .op(n9107) );
  nand4_1 U9280 ( .ip1(n9110), .ip2(n9109), .ip3(n9108), .ip4(n9107), .op(
        n9111) );
  or4_1 U9281 ( .ip1(n9114), .ip2(n9113), .ip3(n9112), .ip4(n9111), .op(n11112) );
  nand2_1 U9282 ( .ip1(n10828), .ip2(n11112), .op(n9179) );
  nand2_1 U9283 ( .ip1(n9690), .ip2(\cache_data[14][75] ), .op(n9118) );
  nand2_1 U9284 ( .ip1(n9668), .ip2(\cache_data[8][75] ), .op(n9117) );
  nand2_1 U9285 ( .ip1(n9681), .ip2(\cache_data[15][75] ), .op(n9116) );
  nand2_1 U9286 ( .ip1(n9680), .ip2(\cache_data[3][75] ), .op(n9115) );
  nand4_1 U9287 ( .ip1(n9118), .ip2(n9117), .ip3(n9116), .ip4(n9115), .op(
        n9134) );
  nand2_1 U9288 ( .ip1(n9689), .ip2(\cache_data[10][75] ), .op(n9122) );
  nand2_1 U9289 ( .ip1(n9688), .ip2(\cache_data[0][75] ), .op(n9121) );
  nand2_1 U9290 ( .ip1(n8905), .ip2(\cache_data[6][75] ), .op(n9120) );
  nand2_1 U9291 ( .ip1(n9675), .ip2(\cache_data[5][75] ), .op(n9119) );
  nand4_1 U9292 ( .ip1(n9122), .ip2(n9121), .ip3(n9120), .ip4(n9119), .op(
        n9133) );
  nand2_1 U9293 ( .ip1(n12120), .ip2(\cache_data[1][75] ), .op(n9126) );
  nand2_1 U9294 ( .ip1(n9560), .ip2(\cache_data[12][75] ), .op(n9125) );
  nand2_1 U9295 ( .ip1(n9682), .ip2(\cache_data[9][75] ), .op(n9124) );
  nand2_1 U9296 ( .ip1(n9670), .ip2(\cache_data[7][75] ), .op(n9123) );
  nand4_1 U9297 ( .ip1(n9126), .ip2(n9125), .ip3(n9124), .ip4(n9123), .op(
        n9132) );
  nand2_1 U9298 ( .ip1(n9687), .ip2(\cache_data[2][75] ), .op(n9130) );
  nand2_1 U9299 ( .ip1(n11927), .ip2(\cache_data[11][75] ), .op(n9129) );
  nand2_1 U9300 ( .ip1(n12165), .ip2(\cache_data[13][75] ), .op(n9128) );
  nand2_1 U9301 ( .ip1(n12164), .ip2(\cache_data[4][75] ), .op(n9127) );
  nand4_1 U9302 ( .ip1(n9130), .ip2(n9129), .ip3(n9128), .ip4(n9127), .op(
        n9131) );
  nor4_1 U9303 ( .ip1(n9134), .ip2(n9133), .ip3(n9132), .ip4(n9131), .op(
        n11114) );
  nor2_1 U9304 ( .ip1(n11114), .ip2(n10849), .op(n9156) );
  nand2_1 U9305 ( .ip1(n9680), .ip2(\cache_data[3][43] ), .op(n9138) );
  nand2_1 U9306 ( .ip1(n12120), .ip2(\cache_data[1][43] ), .op(n9137) );
  nand2_1 U9307 ( .ip1(n12201), .ip2(\cache_data[4][43] ), .op(n9136) );
  nand2_1 U9308 ( .ip1(n8905), .ip2(\cache_data[6][43] ), .op(n9135) );
  nand4_1 U9309 ( .ip1(n9138), .ip2(n9137), .ip3(n9136), .ip4(n9135), .op(
        n9154) );
  nand2_1 U9310 ( .ip1(n9670), .ip2(\cache_data[7][43] ), .op(n9142) );
  nand2_1 U9311 ( .ip1(n9689), .ip2(\cache_data[10][43] ), .op(n9141) );
  nand2_1 U9312 ( .ip1(n9668), .ip2(\cache_data[8][43] ), .op(n9140) );
  nand2_1 U9313 ( .ip1(n9681), .ip2(\cache_data[15][43] ), .op(n9139) );
  nand4_1 U9314 ( .ip1(n9142), .ip2(n9141), .ip3(n9140), .ip4(n9139), .op(
        n9153) );
  nand2_1 U9315 ( .ip1(n9690), .ip2(\cache_data[14][43] ), .op(n9146) );
  nand2_1 U9316 ( .ip1(n12165), .ip2(\cache_data[13][43] ), .op(n9145) );
  nand2_1 U9317 ( .ip1(n9687), .ip2(\cache_data[2][43] ), .op(n9144) );
  nand2_1 U9318 ( .ip1(n9682), .ip2(\cache_data[9][43] ), .op(n9143) );
  nand4_1 U9319 ( .ip1(n9146), .ip2(n9145), .ip3(n9144), .ip4(n9143), .op(
        n9152) );
  nand2_1 U9320 ( .ip1(n9688), .ip2(\cache_data[0][43] ), .op(n9150) );
  nand2_1 U9321 ( .ip1(n11927), .ip2(\cache_data[11][43] ), .op(n9149) );
  nand2_1 U9322 ( .ip1(n9560), .ip2(\cache_data[12][43] ), .op(n9148) );
  nand2_1 U9323 ( .ip1(n9675), .ip2(\cache_data[5][43] ), .op(n9147) );
  nand4_1 U9324 ( .ip1(n9150), .ip2(n9149), .ip3(n9148), .ip4(n9147), .op(
        n9151) );
  nor4_1 U9325 ( .ip1(n9154), .ip2(n9153), .ip3(n9152), .ip4(n9151), .op(
        n11113) );
  nor2_1 U9326 ( .ip1(n11113), .ip2(n10870), .op(n9155) );
  not_ab_or_c_or_d U9327 ( .ip1(data_wr_mem[11]), .ip2(n10873), .ip3(n9156), 
        .ip4(n9155), .op(n9178) );
  nand2_1 U9328 ( .ip1(n9690), .ip2(\cache_data[14][107] ), .op(n9160) );
  nand2_1 U9329 ( .ip1(n9688), .ip2(\cache_data[0][107] ), .op(n9159) );
  nand2_1 U9330 ( .ip1(n9560), .ip2(\cache_data[12][107] ), .op(n9158) );
  nand2_1 U9331 ( .ip1(n9687), .ip2(\cache_data[2][107] ), .op(n9157) );
  nand4_1 U9332 ( .ip1(n9160), .ip2(n9159), .ip3(n9158), .ip4(n9157), .op(
        n9176) );
  nand2_1 U9333 ( .ip1(n9682), .ip2(\cache_data[9][107] ), .op(n9164) );
  nand2_1 U9334 ( .ip1(n11927), .ip2(\cache_data[11][107] ), .op(n9163) );
  nand2_1 U9335 ( .ip1(n12165), .ip2(\cache_data[13][107] ), .op(n9162) );
  nand2_1 U9336 ( .ip1(n9681), .ip2(\cache_data[15][107] ), .op(n9161) );
  nand4_1 U9337 ( .ip1(n9164), .ip2(n9163), .ip3(n9162), .ip4(n9161), .op(
        n9175) );
  nand2_1 U9338 ( .ip1(n9675), .ip2(\cache_data[5][107] ), .op(n9168) );
  nand2_1 U9339 ( .ip1(n9689), .ip2(\cache_data[10][107] ), .op(n9167) );
  nand2_1 U9340 ( .ip1(n9680), .ip2(\cache_data[3][107] ), .op(n9166) );
  nand2_1 U9341 ( .ip1(n12120), .ip2(\cache_data[1][107] ), .op(n9165) );
  nand4_1 U9342 ( .ip1(n9168), .ip2(n9167), .ip3(n9166), .ip4(n9165), .op(
        n9174) );
  nand2_1 U9343 ( .ip1(n9668), .ip2(\cache_data[8][107] ), .op(n9172) );
  nand2_1 U9344 ( .ip1(n12201), .ip2(\cache_data[4][107] ), .op(n9171) );
  nand2_1 U9345 ( .ip1(n10305), .ip2(\cache_data[6][107] ), .op(n9170) );
  nand2_1 U9346 ( .ip1(n9670), .ip2(\cache_data[7][107] ), .op(n9169) );
  nand4_1 U9347 ( .ip1(n9172), .ip2(n9171), .ip3(n9170), .ip4(n9169), .op(
        n9173) );
  or4_1 U9348 ( .ip1(n9176), .ip2(n9175), .ip3(n9174), .ip4(n9173), .op(n11117) );
  nand2_1 U9349 ( .ip1(n10894), .ip2(n11117), .op(n9177) );
  nand3_1 U9350 ( .ip1(n9179), .ip2(n9178), .ip3(n9177), .op(n7437) );
  nand2_1 U9351 ( .ip1(data_wr_mem[12]), .ip2(n10873), .op(n9264) );
  nand2_1 U9352 ( .ip1(n9690), .ip2(\cache_data[14][108] ), .op(n9183) );
  nand2_1 U9353 ( .ip1(n9688), .ip2(\cache_data[0][108] ), .op(n9182) );
  nand2_1 U9354 ( .ip1(n12179), .ip2(\cache_data[6][108] ), .op(n9181) );
  nand2_1 U9355 ( .ip1(n9682), .ip2(\cache_data[9][108] ), .op(n9180) );
  nand4_1 U9356 ( .ip1(n9183), .ip2(n9182), .ip3(n9181), .ip4(n9180), .op(
        n9199) );
  nand2_1 U9357 ( .ip1(n9681), .ip2(\cache_data[15][108] ), .op(n9187) );
  nand2_1 U9358 ( .ip1(n9668), .ip2(\cache_data[8][108] ), .op(n9186) );
  nand2_1 U9359 ( .ip1(n9675), .ip2(\cache_data[5][108] ), .op(n9185) );
  nand2_1 U9360 ( .ip1(n12243), .ip2(\cache_data[4][108] ), .op(n9184) );
  nand4_1 U9361 ( .ip1(n9187), .ip2(n9186), .ip3(n9185), .ip4(n9184), .op(
        n9198) );
  nand2_1 U9362 ( .ip1(n9680), .ip2(\cache_data[3][108] ), .op(n9191) );
  nand2_1 U9363 ( .ip1(n12227), .ip2(\cache_data[12][108] ), .op(n9190) );
  nand2_1 U9364 ( .ip1(n9687), .ip2(\cache_data[2][108] ), .op(n9189) );
  nand2_1 U9365 ( .ip1(n9689), .ip2(\cache_data[10][108] ), .op(n9188) );
  nand4_1 U9366 ( .ip1(n9191), .ip2(n9190), .ip3(n9189), .ip4(n9188), .op(
        n9197) );
  nand2_1 U9367 ( .ip1(n12142), .ip2(\cache_data[13][108] ), .op(n9195) );
  nand2_1 U9368 ( .ip1(n11927), .ip2(\cache_data[11][108] ), .op(n9194) );
  nand2_1 U9369 ( .ip1(n12120), .ip2(\cache_data[1][108] ), .op(n9193) );
  nand2_1 U9370 ( .ip1(n9670), .ip2(\cache_data[7][108] ), .op(n9192) );
  nand4_1 U9371 ( .ip1(n9195), .ip2(n9194), .ip3(n9193), .ip4(n9192), .op(
        n9196) );
  or4_1 U9372 ( .ip1(n9199), .ip2(n9198), .ip3(n9197), .ip4(n9196), .op(n11121) );
  nand2_1 U9373 ( .ip1(n9682), .ip2(\cache_data[9][76] ), .op(n9203) );
  nand2_1 U9374 ( .ip1(n12227), .ip2(\cache_data[12][76] ), .op(n9202) );
  nand2_1 U9375 ( .ip1(n9670), .ip2(\cache_data[7][76] ), .op(n9201) );
  nand2_1 U9376 ( .ip1(n12201), .ip2(\cache_data[4][76] ), .op(n9200) );
  nand4_1 U9377 ( .ip1(n9203), .ip2(n9202), .ip3(n9201), .ip4(n9200), .op(
        n9219) );
  nand2_1 U9378 ( .ip1(n12179), .ip2(\cache_data[6][76] ), .op(n9207) );
  nand2_1 U9379 ( .ip1(n9687), .ip2(\cache_data[2][76] ), .op(n9206) );
  nand2_1 U9380 ( .ip1(n9689), .ip2(\cache_data[10][76] ), .op(n9205) );
  nand2_1 U9381 ( .ip1(n9680), .ip2(\cache_data[3][76] ), .op(n9204) );
  nand4_1 U9382 ( .ip1(n9207), .ip2(n9206), .ip3(n9205), .ip4(n9204), .op(
        n9218) );
  nand2_1 U9383 ( .ip1(n11927), .ip2(\cache_data[11][76] ), .op(n9211) );
  nand2_1 U9384 ( .ip1(n9681), .ip2(\cache_data[15][76] ), .op(n9210) );
  nand2_1 U9385 ( .ip1(n12142), .ip2(\cache_data[13][76] ), .op(n9209) );
  nand2_1 U9386 ( .ip1(n9690), .ip2(\cache_data[14][76] ), .op(n9208) );
  nand4_1 U9387 ( .ip1(n9211), .ip2(n9210), .ip3(n9209), .ip4(n9208), .op(
        n9217) );
  nand2_1 U9388 ( .ip1(n9668), .ip2(\cache_data[8][76] ), .op(n9215) );
  nand2_1 U9389 ( .ip1(n12120), .ip2(\cache_data[1][76] ), .op(n9214) );
  nand2_1 U9390 ( .ip1(n9675), .ip2(\cache_data[5][76] ), .op(n9213) );
  nand2_1 U9391 ( .ip1(n9688), .ip2(\cache_data[0][76] ), .op(n9212) );
  nand4_1 U9392 ( .ip1(n9215), .ip2(n9214), .ip3(n9213), .ip4(n9212), .op(
        n9216) );
  nor4_1 U9393 ( .ip1(n9219), .ip2(n9218), .ip3(n9217), .ip4(n9216), .op(
        n11122) );
  nor2_1 U9394 ( .ip1(n11122), .ip2(n10849), .op(n9241) );
  nand2_1 U9395 ( .ip1(n9689), .ip2(\cache_data[10][44] ), .op(n9223) );
  nand2_1 U9396 ( .ip1(n9680), .ip2(\cache_data[3][44] ), .op(n9222) );
  nand2_1 U9397 ( .ip1(n9681), .ip2(\cache_data[15][44] ), .op(n9221) );
  nand2_1 U9398 ( .ip1(n12201), .ip2(\cache_data[4][44] ), .op(n9220) );
  nand4_1 U9399 ( .ip1(n9223), .ip2(n9222), .ip3(n9221), .ip4(n9220), .op(
        n9239) );
  nand2_1 U9400 ( .ip1(n9687), .ip2(\cache_data[2][44] ), .op(n9227) );
  inv_1 U9401 ( .ip(n8151), .op(n9669) );
  nand2_1 U9402 ( .ip1(n9669), .ip2(\cache_data[11][44] ), .op(n9226) );
  nand2_1 U9403 ( .ip1(n12165), .ip2(\cache_data[13][44] ), .op(n9225) );
  nand2_1 U9404 ( .ip1(n9682), .ip2(\cache_data[9][44] ), .op(n9224) );
  nand4_1 U9405 ( .ip1(n9227), .ip2(n9226), .ip3(n9225), .ip4(n9224), .op(
        n9238) );
  nand2_1 U9406 ( .ip1(n12227), .ip2(\cache_data[12][44] ), .op(n9231) );
  nand2_1 U9407 ( .ip1(n12120), .ip2(\cache_data[1][44] ), .op(n9230) );
  nand2_1 U9408 ( .ip1(n9670), .ip2(\cache_data[7][44] ), .op(n9229) );
  nand2_1 U9409 ( .ip1(n9668), .ip2(\cache_data[8][44] ), .op(n9228) );
  nand4_1 U9410 ( .ip1(n9231), .ip2(n9230), .ip3(n9229), .ip4(n9228), .op(
        n9237) );
  nand2_1 U9411 ( .ip1(n9688), .ip2(\cache_data[0][44] ), .op(n9235) );
  nand2_1 U9412 ( .ip1(n12179), .ip2(\cache_data[6][44] ), .op(n9234) );
  nand2_1 U9413 ( .ip1(n9690), .ip2(\cache_data[14][44] ), .op(n9233) );
  nand2_1 U9414 ( .ip1(n9675), .ip2(\cache_data[5][44] ), .op(n9232) );
  nand4_1 U9415 ( .ip1(n9235), .ip2(n9234), .ip3(n9233), .ip4(n9232), .op(
        n9236) );
  nor4_1 U9416 ( .ip1(n9239), .ip2(n9238), .ip3(n9237), .ip4(n9236), .op(
        n11123) );
  nor2_1 U9417 ( .ip1(n11123), .ip2(n10870), .op(n9240) );
  not_ab_or_c_or_d U9418 ( .ip1(n10894), .ip2(n11121), .ip3(n9241), .ip4(n9240), .op(n9263) );
  nand2_1 U9419 ( .ip1(n12096), .ip2(\cache_data[11][12] ), .op(n9245) );
  nand2_1 U9420 ( .ip1(n9680), .ip2(\cache_data[3][12] ), .op(n9244) );
  nand2_1 U9421 ( .ip1(n12207), .ip2(\cache_data[12][12] ), .op(n9243) );
  nand2_1 U9422 ( .ip1(n12179), .ip2(\cache_data[6][12] ), .op(n9242) );
  nand4_1 U9423 ( .ip1(n9245), .ip2(n9244), .ip3(n9243), .ip4(n9242), .op(
        n9261) );
  nand2_1 U9424 ( .ip1(n9687), .ip2(\cache_data[2][12] ), .op(n9249) );
  nand2_1 U9425 ( .ip1(n9682), .ip2(\cache_data[9][12] ), .op(n9248) );
  nand2_1 U9426 ( .ip1(n9690), .ip2(\cache_data[14][12] ), .op(n9247) );
  nand2_1 U9427 ( .ip1(n9675), .ip2(\cache_data[5][12] ), .op(n9246) );
  nand4_1 U9428 ( .ip1(n9249), .ip2(n9248), .ip3(n9247), .ip4(n9246), .op(
        n9260) );
  nand2_1 U9429 ( .ip1(n12201), .ip2(\cache_data[4][12] ), .op(n9253) );
  nand2_1 U9430 ( .ip1(n9688), .ip2(\cache_data[0][12] ), .op(n9252) );
  nand2_1 U9431 ( .ip1(n9689), .ip2(\cache_data[10][12] ), .op(n9251) );
  nand2_1 U9432 ( .ip1(n9681), .ip2(\cache_data[15][12] ), .op(n9250) );
  nand4_1 U9433 ( .ip1(n9253), .ip2(n9252), .ip3(n9251), .ip4(n9250), .op(
        n9259) );
  nand2_1 U9434 ( .ip1(n12142), .ip2(\cache_data[13][12] ), .op(n9257) );
  nand2_1 U9435 ( .ip1(n9670), .ip2(\cache_data[7][12] ), .op(n9256) );
  nand2_1 U9436 ( .ip1(n9668), .ip2(\cache_data[8][12] ), .op(n9255) );
  nand2_1 U9437 ( .ip1(n12120), .ip2(\cache_data[1][12] ), .op(n9254) );
  nand4_1 U9438 ( .ip1(n9257), .ip2(n9256), .ip3(n9255), .ip4(n9254), .op(
        n9258) );
  or4_1 U9439 ( .ip1(n9261), .ip2(n9260), .ip3(n9259), .ip4(n9258), .op(n11126) );
  nand2_1 U9440 ( .ip1(n10828), .ip2(n11126), .op(n9262) );
  nand3_1 U9441 ( .ip1(n9264), .ip2(n9263), .ip3(n9262), .op(n7436) );
  nand2_1 U9442 ( .ip1(n9689), .ip2(\cache_data[10][13] ), .op(n9268) );
  nand2_1 U9443 ( .ip1(n9681), .ip2(\cache_data[15][13] ), .op(n9267) );
  nand2_1 U9444 ( .ip1(n9675), .ip2(\cache_data[5][13] ), .op(n9266) );
  nand2_1 U9445 ( .ip1(n9670), .ip2(\cache_data[7][13] ), .op(n9265) );
  nand4_1 U9446 ( .ip1(n9268), .ip2(n9267), .ip3(n9266), .ip4(n9265), .op(
        n9284) );
  nand2_1 U9447 ( .ip1(n9687), .ip2(\cache_data[2][13] ), .op(n9272) );
  nand2_1 U9448 ( .ip1(n12179), .ip2(\cache_data[6][13] ), .op(n9271) );
  nand2_1 U9449 ( .ip1(n12201), .ip2(\cache_data[4][13] ), .op(n9270) );
  nand2_1 U9450 ( .ip1(n9688), .ip2(\cache_data[0][13] ), .op(n9269) );
  nand4_1 U9451 ( .ip1(n9272), .ip2(n9271), .ip3(n9270), .ip4(n9269), .op(
        n9283) );
  nand2_1 U9452 ( .ip1(n9690), .ip2(\cache_data[14][13] ), .op(n9276) );
  nand2_1 U9453 ( .ip1(n12096), .ip2(\cache_data[11][13] ), .op(n9275) );
  nand2_1 U9454 ( .ip1(n12120), .ip2(\cache_data[1][13] ), .op(n9274) );
  nand2_1 U9455 ( .ip1(n9668), .ip2(\cache_data[8][13] ), .op(n9273) );
  nand4_1 U9456 ( .ip1(n9276), .ip2(n9275), .ip3(n9274), .ip4(n9273), .op(
        n9282) );
  nand2_1 U9457 ( .ip1(n12142), .ip2(\cache_data[13][13] ), .op(n9280) );
  nand2_1 U9458 ( .ip1(n12207), .ip2(\cache_data[12][13] ), .op(n9279) );
  nand2_1 U9459 ( .ip1(n9680), .ip2(\cache_data[3][13] ), .op(n9278) );
  nand2_1 U9460 ( .ip1(n9682), .ip2(\cache_data[9][13] ), .op(n9277) );
  nand4_1 U9461 ( .ip1(n9280), .ip2(n9279), .ip3(n9278), .ip4(n9277), .op(
        n9281) );
  or4_1 U9462 ( .ip1(n9284), .ip2(n9283), .ip3(n9282), .ip4(n9281), .op(n11130) );
  nand2_1 U9463 ( .ip1(n10828), .ip2(n11130), .op(n9349) );
  nand2_1 U9464 ( .ip1(n12120), .ip2(\cache_data[1][77] ), .op(n9288) );
  nand2_1 U9465 ( .ip1(n9670), .ip2(\cache_data[7][77] ), .op(n9287) );
  nand2_1 U9466 ( .ip1(n9682), .ip2(\cache_data[9][77] ), .op(n9286) );
  nand2_1 U9467 ( .ip1(n9681), .ip2(\cache_data[15][77] ), .op(n9285) );
  nand4_1 U9468 ( .ip1(n9288), .ip2(n9287), .ip3(n9286), .ip4(n9285), .op(
        n9304) );
  nand2_1 U9469 ( .ip1(n9669), .ip2(\cache_data[11][77] ), .op(n9292) );
  nand2_1 U9470 ( .ip1(n9688), .ip2(\cache_data[0][77] ), .op(n9291) );
  nand2_1 U9471 ( .ip1(n8905), .ip2(\cache_data[6][77] ), .op(n9290) );
  nand2_1 U9472 ( .ip1(n9689), .ip2(\cache_data[10][77] ), .op(n9289) );
  nand4_1 U9473 ( .ip1(n9292), .ip2(n9291), .ip3(n9290), .ip4(n9289), .op(
        n9303) );
  nand2_1 U9474 ( .ip1(n9680), .ip2(\cache_data[3][77] ), .op(n9296) );
  nand2_1 U9475 ( .ip1(n9675), .ip2(\cache_data[5][77] ), .op(n9295) );
  nand2_1 U9476 ( .ip1(n9690), .ip2(\cache_data[14][77] ), .op(n9294) );
  nand2_1 U9477 ( .ip1(n9668), .ip2(\cache_data[8][77] ), .op(n9293) );
  nand4_1 U9478 ( .ip1(n9296), .ip2(n9295), .ip3(n9294), .ip4(n9293), .op(
        n9302) );
  nand2_1 U9479 ( .ip1(n9687), .ip2(\cache_data[2][77] ), .op(n9300) );
  nand2_1 U9480 ( .ip1(n12243), .ip2(\cache_data[4][77] ), .op(n9299) );
  nand2_1 U9481 ( .ip1(n12227), .ip2(\cache_data[12][77] ), .op(n9298) );
  nand2_1 U9482 ( .ip1(n12142), .ip2(\cache_data[13][77] ), .op(n9297) );
  nand4_1 U9483 ( .ip1(n9300), .ip2(n9299), .ip3(n9298), .ip4(n9297), .op(
        n9301) );
  nor4_1 U9484 ( .ip1(n9304), .ip2(n9303), .ip3(n9302), .ip4(n9301), .op(
        n11131) );
  nor2_1 U9485 ( .ip1(n11131), .ip2(n10849), .op(n9326) );
  nand2_1 U9486 ( .ip1(n8905), .ip2(\cache_data[6][45] ), .op(n9308) );
  nand2_1 U9487 ( .ip1(n9688), .ip2(\cache_data[0][45] ), .op(n9307) );
  nand2_1 U9488 ( .ip1(n9689), .ip2(\cache_data[10][45] ), .op(n9306) );
  nand2_1 U9489 ( .ip1(n9668), .ip2(\cache_data[8][45] ), .op(n9305) );
  nand4_1 U9490 ( .ip1(n9308), .ip2(n9307), .ip3(n9306), .ip4(n9305), .op(
        n9324) );
  nand2_1 U9491 ( .ip1(n11927), .ip2(\cache_data[11][45] ), .op(n9312) );
  nand2_1 U9492 ( .ip1(n9680), .ip2(\cache_data[3][45] ), .op(n9311) );
  nand2_1 U9493 ( .ip1(n9681), .ip2(\cache_data[15][45] ), .op(n9310) );
  nand2_1 U9494 ( .ip1(n9687), .ip2(\cache_data[2][45] ), .op(n9309) );
  nand4_1 U9495 ( .ip1(n9312), .ip2(n9311), .ip3(n9310), .ip4(n9309), .op(
        n9323) );
  nand2_1 U9496 ( .ip1(n12243), .ip2(\cache_data[4][45] ), .op(n9316) );
  nand2_1 U9497 ( .ip1(n12227), .ip2(\cache_data[12][45] ), .op(n9315) );
  nand2_1 U9498 ( .ip1(n12120), .ip2(\cache_data[1][45] ), .op(n9314) );
  nand2_1 U9499 ( .ip1(n9682), .ip2(\cache_data[9][45] ), .op(n9313) );
  nand4_1 U9500 ( .ip1(n9316), .ip2(n9315), .ip3(n9314), .ip4(n9313), .op(
        n9322) );
  nand2_1 U9501 ( .ip1(n12142), .ip2(\cache_data[13][45] ), .op(n9320) );
  nand2_1 U9502 ( .ip1(n9670), .ip2(\cache_data[7][45] ), .op(n9319) );
  nand2_1 U9503 ( .ip1(n9690), .ip2(\cache_data[14][45] ), .op(n9318) );
  nand2_1 U9504 ( .ip1(n9675), .ip2(\cache_data[5][45] ), .op(n9317) );
  nand4_1 U9505 ( .ip1(n9320), .ip2(n9319), .ip3(n9318), .ip4(n9317), .op(
        n9321) );
  nor4_1 U9506 ( .ip1(n9324), .ip2(n9323), .ip3(n9322), .ip4(n9321), .op(
        n11132) );
  nor2_1 U9507 ( .ip1(n11132), .ip2(n10870), .op(n9325) );
  not_ab_or_c_or_d U9508 ( .ip1(data_wr_mem[13]), .ip2(n10873), .ip3(n9326), 
        .ip4(n9325), .op(n9348) );
  nand2_1 U9509 ( .ip1(n9668), .ip2(\cache_data[8][109] ), .op(n9330) );
  nand2_1 U9510 ( .ip1(n9690), .ip2(\cache_data[14][109] ), .op(n9329) );
  nand2_1 U9511 ( .ip1(n9680), .ip2(\cache_data[3][109] ), .op(n9328) );
  nand2_1 U9512 ( .ip1(n12227), .ip2(\cache_data[12][109] ), .op(n9327) );
  nand4_1 U9513 ( .ip1(n9330), .ip2(n9329), .ip3(n9328), .ip4(n9327), .op(
        n9346) );
  nand2_1 U9514 ( .ip1(n9688), .ip2(\cache_data[0][109] ), .op(n9334) );
  nand2_1 U9515 ( .ip1(n9681), .ip2(\cache_data[15][109] ), .op(n9333) );
  nand2_1 U9516 ( .ip1(n9689), .ip2(\cache_data[10][109] ), .op(n9332) );
  nand2_1 U9517 ( .ip1(n9687), .ip2(\cache_data[2][109] ), .op(n9331) );
  nand4_1 U9518 ( .ip1(n9334), .ip2(n9333), .ip3(n9332), .ip4(n9331), .op(
        n9345) );
  nand2_1 U9519 ( .ip1(n12120), .ip2(\cache_data[1][109] ), .op(n9338) );
  nand2_1 U9520 ( .ip1(n9670), .ip2(\cache_data[7][109] ), .op(n9337) );
  nand2_1 U9521 ( .ip1(n9682), .ip2(\cache_data[9][109] ), .op(n9336) );
  nand2_1 U9522 ( .ip1(n11927), .ip2(\cache_data[11][109] ), .op(n9335) );
  nand4_1 U9523 ( .ip1(n9338), .ip2(n9337), .ip3(n9336), .ip4(n9335), .op(
        n9344) );
  nand2_1 U9524 ( .ip1(n12142), .ip2(\cache_data[13][109] ), .op(n9342) );
  nand2_1 U9525 ( .ip1(n12179), .ip2(\cache_data[6][109] ), .op(n9341) );
  nand2_1 U9526 ( .ip1(n12243), .ip2(\cache_data[4][109] ), .op(n9340) );
  nand2_1 U9527 ( .ip1(n9675), .ip2(\cache_data[5][109] ), .op(n9339) );
  nand4_1 U9528 ( .ip1(n9342), .ip2(n9341), .ip3(n9340), .ip4(n9339), .op(
        n9343) );
  or4_1 U9529 ( .ip1(n9346), .ip2(n9345), .ip3(n9344), .ip4(n9343), .op(n11135) );
  nand2_1 U9530 ( .ip1(n10894), .ip2(n11135), .op(n9347) );
  nand3_1 U9531 ( .ip1(n9349), .ip2(n9348), .ip3(n9347), .op(n7435) );
  nand2_1 U9532 ( .ip1(data_wr_mem[14]), .ip2(n10873), .op(n9434) );
  nand2_1 U9533 ( .ip1(n12120), .ip2(\cache_data[1][14] ), .op(n9353) );
  nand2_1 U9534 ( .ip1(n9682), .ip2(\cache_data[9][14] ), .op(n9352) );
  nand2_1 U9535 ( .ip1(n12227), .ip2(\cache_data[12][14] ), .op(n9351) );
  nand2_1 U9536 ( .ip1(n9690), .ip2(\cache_data[14][14] ), .op(n9350) );
  nand4_1 U9537 ( .ip1(n9353), .ip2(n9352), .ip3(n9351), .ip4(n9350), .op(
        n9369) );
  nand2_1 U9538 ( .ip1(n12179), .ip2(\cache_data[6][14] ), .op(n9357) );
  nand2_1 U9539 ( .ip1(n9675), .ip2(\cache_data[5][14] ), .op(n9356) );
  nand2_1 U9540 ( .ip1(n12243), .ip2(\cache_data[4][14] ), .op(n9355) );
  nand2_1 U9541 ( .ip1(n9680), .ip2(\cache_data[3][14] ), .op(n9354) );
  nand4_1 U9542 ( .ip1(n9357), .ip2(n9356), .ip3(n9355), .ip4(n9354), .op(
        n9368) );
  nand2_1 U9543 ( .ip1(n11927), .ip2(\cache_data[11][14] ), .op(n9361) );
  nand2_1 U9544 ( .ip1(n9687), .ip2(\cache_data[2][14] ), .op(n9360) );
  nand2_1 U9545 ( .ip1(n9689), .ip2(\cache_data[10][14] ), .op(n9359) );
  nand2_1 U9546 ( .ip1(n9688), .ip2(\cache_data[0][14] ), .op(n9358) );
  nand4_1 U9547 ( .ip1(n9361), .ip2(n9360), .ip3(n9359), .ip4(n9358), .op(
        n9367) );
  nand2_1 U9548 ( .ip1(n9670), .ip2(\cache_data[7][14] ), .op(n9365) );
  nand2_1 U9549 ( .ip1(n9668), .ip2(\cache_data[8][14] ), .op(n9364) );
  nand2_1 U9550 ( .ip1(n9681), .ip2(\cache_data[15][14] ), .op(n9363) );
  nand2_1 U9551 ( .ip1(n12142), .ip2(\cache_data[13][14] ), .op(n9362) );
  nand4_1 U9552 ( .ip1(n9365), .ip2(n9364), .ip3(n9363), .ip4(n9362), .op(
        n9366) );
  or4_1 U9553 ( .ip1(n9369), .ip2(n9368), .ip3(n9367), .ip4(n9366), .op(n11139) );
  nand2_1 U9554 ( .ip1(n9681), .ip2(\cache_data[15][46] ), .op(n9373) );
  nand2_1 U9555 ( .ip1(n9560), .ip2(\cache_data[12][46] ), .op(n9372) );
  nand2_1 U9556 ( .ip1(n12165), .ip2(\cache_data[13][46] ), .op(n9371) );
  nand2_1 U9557 ( .ip1(n12179), .ip2(\cache_data[6][46] ), .op(n9370) );
  nand4_1 U9558 ( .ip1(n9373), .ip2(n9372), .ip3(n9371), .ip4(n9370), .op(
        n9389) );
  nand2_1 U9559 ( .ip1(n9668), .ip2(\cache_data[8][46] ), .op(n9377) );
  nand2_1 U9560 ( .ip1(n9689), .ip2(\cache_data[10][46] ), .op(n9376) );
  nand2_1 U9561 ( .ip1(n9687), .ip2(\cache_data[2][46] ), .op(n9375) );
  nand2_1 U9562 ( .ip1(n11927), .ip2(\cache_data[11][46] ), .op(n9374) );
  nand4_1 U9563 ( .ip1(n9377), .ip2(n9376), .ip3(n9375), .ip4(n9374), .op(
        n9388) );
  nand2_1 U9564 ( .ip1(n12243), .ip2(\cache_data[4][46] ), .op(n9381) );
  nand2_1 U9565 ( .ip1(n9670), .ip2(\cache_data[7][46] ), .op(n9380) );
  nand2_1 U9566 ( .ip1(n9690), .ip2(\cache_data[14][46] ), .op(n9379) );
  nand2_1 U9567 ( .ip1(n9688), .ip2(\cache_data[0][46] ), .op(n9378) );
  nand4_1 U9568 ( .ip1(n9381), .ip2(n9380), .ip3(n9379), .ip4(n9378), .op(
        n9387) );
  nand2_1 U9569 ( .ip1(n9680), .ip2(\cache_data[3][46] ), .op(n9385) );
  nand2_1 U9570 ( .ip1(n9682), .ip2(\cache_data[9][46] ), .op(n9384) );
  nand2_1 U9571 ( .ip1(n9675), .ip2(\cache_data[5][46] ), .op(n9383) );
  nand2_1 U9572 ( .ip1(n12120), .ip2(\cache_data[1][46] ), .op(n9382) );
  nand4_1 U9573 ( .ip1(n9385), .ip2(n9384), .ip3(n9383), .ip4(n9382), .op(
        n9386) );
  nor4_1 U9574 ( .ip1(n9389), .ip2(n9388), .ip3(n9387), .ip4(n9386), .op(
        n11140) );
  nor2_1 U9575 ( .ip1(n11140), .ip2(n10870), .op(n9411) );
  nand2_1 U9576 ( .ip1(n9682), .ip2(\cache_data[9][78] ), .op(n9393) );
  nand2_1 U9577 ( .ip1(n9669), .ip2(\cache_data[11][78] ), .op(n9392) );
  nand2_1 U9578 ( .ip1(n9687), .ip2(\cache_data[2][78] ), .op(n9391) );
  nand2_1 U9579 ( .ip1(n9560), .ip2(\cache_data[12][78] ), .op(n9390) );
  nand4_1 U9580 ( .ip1(n9393), .ip2(n9392), .ip3(n9391), .ip4(n9390), .op(
        n9409) );
  nand2_1 U9581 ( .ip1(n9689), .ip2(\cache_data[10][78] ), .op(n9397) );
  nand2_1 U9582 ( .ip1(n9668), .ip2(\cache_data[8][78] ), .op(n9396) );
  nand2_1 U9583 ( .ip1(n12120), .ip2(\cache_data[1][78] ), .op(n9395) );
  nand2_1 U9584 ( .ip1(n12243), .ip2(\cache_data[4][78] ), .op(n9394) );
  nand4_1 U9585 ( .ip1(n9397), .ip2(n9396), .ip3(n9395), .ip4(n9394), .op(
        n9408) );
  nand2_1 U9586 ( .ip1(n9680), .ip2(\cache_data[3][78] ), .op(n9401) );
  nand2_1 U9587 ( .ip1(n12142), .ip2(\cache_data[13][78] ), .op(n9400) );
  nand2_1 U9588 ( .ip1(n9675), .ip2(\cache_data[5][78] ), .op(n9399) );
  nand2_1 U9589 ( .ip1(n9690), .ip2(\cache_data[14][78] ), .op(n9398) );
  nand4_1 U9590 ( .ip1(n9401), .ip2(n9400), .ip3(n9399), .ip4(n9398), .op(
        n9407) );
  nand2_1 U9591 ( .ip1(n12179), .ip2(\cache_data[6][78] ), .op(n9405) );
  nand2_1 U9592 ( .ip1(n9688), .ip2(\cache_data[0][78] ), .op(n9404) );
  nand2_1 U9593 ( .ip1(n9681), .ip2(\cache_data[15][78] ), .op(n9403) );
  nand2_1 U9594 ( .ip1(n9670), .ip2(\cache_data[7][78] ), .op(n9402) );
  nand4_1 U9595 ( .ip1(n9405), .ip2(n9404), .ip3(n9403), .ip4(n9402), .op(
        n9406) );
  nor4_1 U9596 ( .ip1(n9409), .ip2(n9408), .ip3(n9407), .ip4(n9406), .op(
        n11141) );
  nor2_1 U9597 ( .ip1(n11141), .ip2(n10849), .op(n9410) );
  not_ab_or_c_or_d U9598 ( .ip1(n10828), .ip2(n11139), .ip3(n9411), .ip4(n9410), .op(n9433) );
  nand2_1 U9599 ( .ip1(n11927), .ip2(\cache_data[11][110] ), .op(n9415) );
  nand2_1 U9600 ( .ip1(n9680), .ip2(\cache_data[3][110] ), .op(n9414) );
  nand2_1 U9601 ( .ip1(n9688), .ip2(\cache_data[0][110] ), .op(n9413) );
  nand2_1 U9602 ( .ip1(n9690), .ip2(\cache_data[14][110] ), .op(n9412) );
  nand4_1 U9603 ( .ip1(n9415), .ip2(n9414), .ip3(n9413), .ip4(n9412), .op(
        n9431) );
  nand2_1 U9604 ( .ip1(n9675), .ip2(\cache_data[5][110] ), .op(n9419) );
  nand2_1 U9605 ( .ip1(n9670), .ip2(\cache_data[7][110] ), .op(n9418) );
  nand2_1 U9606 ( .ip1(n12243), .ip2(\cache_data[4][110] ), .op(n9417) );
  nand2_1 U9607 ( .ip1(n12142), .ip2(\cache_data[13][110] ), .op(n9416) );
  nand4_1 U9608 ( .ip1(n9419), .ip2(n9418), .ip3(n9417), .ip4(n9416), .op(
        n9430) );
  nand2_1 U9609 ( .ip1(n12227), .ip2(\cache_data[12][110] ), .op(n9423) );
  nand2_1 U9610 ( .ip1(n12179), .ip2(\cache_data[6][110] ), .op(n9422) );
  nand2_1 U9611 ( .ip1(n9668), .ip2(\cache_data[8][110] ), .op(n9421) );
  nand2_1 U9612 ( .ip1(n9687), .ip2(\cache_data[2][110] ), .op(n9420) );
  nand4_1 U9613 ( .ip1(n9423), .ip2(n9422), .ip3(n9421), .ip4(n9420), .op(
        n9429) );
  nand2_1 U9614 ( .ip1(n12120), .ip2(\cache_data[1][110] ), .op(n9427) );
  nand2_1 U9615 ( .ip1(n9682), .ip2(\cache_data[9][110] ), .op(n9426) );
  nand2_1 U9616 ( .ip1(n9689), .ip2(\cache_data[10][110] ), .op(n9425) );
  nand2_1 U9617 ( .ip1(n9681), .ip2(\cache_data[15][110] ), .op(n9424) );
  nand4_1 U9618 ( .ip1(n9427), .ip2(n9426), .ip3(n9425), .ip4(n9424), .op(
        n9428) );
  or4_1 U9619 ( .ip1(n9431), .ip2(n9430), .ip3(n9429), .ip4(n9428), .op(n11144) );
  nand2_1 U9620 ( .ip1(n10894), .ip2(n11144), .op(n9432) );
  nand3_1 U9621 ( .ip1(n9434), .ip2(n9433), .ip3(n9432), .op(n7434) );
  nand2_1 U9622 ( .ip1(n12120), .ip2(\cache_data[1][15] ), .op(n9438) );
  nand2_1 U9623 ( .ip1(n9688), .ip2(\cache_data[0][15] ), .op(n9437) );
  nand2_1 U9624 ( .ip1(n9668), .ip2(\cache_data[8][15] ), .op(n9436) );
  nand2_1 U9625 ( .ip1(n9669), .ip2(\cache_data[11][15] ), .op(n9435) );
  nand4_1 U9626 ( .ip1(n9438), .ip2(n9437), .ip3(n9436), .ip4(n9435), .op(
        n9454) );
  nand2_1 U9627 ( .ip1(n12179), .ip2(\cache_data[6][15] ), .op(n9442) );
  nand2_1 U9628 ( .ip1(n9689), .ip2(\cache_data[10][15] ), .op(n9441) );
  nand2_1 U9629 ( .ip1(n12207), .ip2(\cache_data[12][15] ), .op(n9440) );
  nand2_1 U9630 ( .ip1(n9687), .ip2(\cache_data[2][15] ), .op(n9439) );
  nand4_1 U9631 ( .ip1(n9442), .ip2(n9441), .ip3(n9440), .ip4(n9439), .op(
        n9453) );
  nand2_1 U9632 ( .ip1(n9675), .ip2(\cache_data[5][15] ), .op(n9446) );
  nand2_1 U9633 ( .ip1(n9670), .ip2(\cache_data[7][15] ), .op(n9445) );
  nand2_1 U9634 ( .ip1(n9690), .ip2(\cache_data[14][15] ), .op(n9444) );
  nand2_1 U9635 ( .ip1(n9682), .ip2(\cache_data[9][15] ), .op(n9443) );
  nand4_1 U9636 ( .ip1(n9446), .ip2(n9445), .ip3(n9444), .ip4(n9443), .op(
        n9452) );
  nand2_1 U9637 ( .ip1(n12142), .ip2(\cache_data[13][15] ), .op(n9450) );
  nand2_1 U9638 ( .ip1(n9680), .ip2(\cache_data[3][15] ), .op(n9449) );
  nand2_1 U9639 ( .ip1(n9681), .ip2(\cache_data[15][15] ), .op(n9448) );
  nand2_1 U9640 ( .ip1(n12201), .ip2(\cache_data[4][15] ), .op(n9447) );
  nand4_1 U9641 ( .ip1(n9450), .ip2(n9449), .ip3(n9448), .ip4(n9447), .op(
        n9451) );
  or4_1 U9642 ( .ip1(n9454), .ip2(n9453), .ip3(n9452), .ip4(n9451), .op(n11148) );
  nand2_1 U9643 ( .ip1(n10828), .ip2(n11148), .op(n9519) );
  nand2_1 U9644 ( .ip1(n12227), .ip2(\cache_data[12][79] ), .op(n9458) );
  nand2_1 U9645 ( .ip1(n9669), .ip2(\cache_data[11][79] ), .op(n9457) );
  nand2_1 U9646 ( .ip1(n9668), .ip2(\cache_data[8][79] ), .op(n9456) );
  nand2_1 U9647 ( .ip1(n9687), .ip2(\cache_data[2][79] ), .op(n9455) );
  nand4_1 U9648 ( .ip1(n9458), .ip2(n9457), .ip3(n9456), .ip4(n9455), .op(
        n9474) );
  nand2_1 U9649 ( .ip1(n9675), .ip2(\cache_data[5][79] ), .op(n9462) );
  nand2_1 U9650 ( .ip1(n9670), .ip2(\cache_data[7][79] ), .op(n9461) );
  nand2_1 U9651 ( .ip1(n12120), .ip2(\cache_data[1][79] ), .op(n9460) );
  nand2_1 U9652 ( .ip1(n9680), .ip2(\cache_data[3][79] ), .op(n9459) );
  nand4_1 U9653 ( .ip1(n9462), .ip2(n9461), .ip3(n9460), .ip4(n9459), .op(
        n9473) );
  nand2_1 U9654 ( .ip1(n12179), .ip2(\cache_data[6][79] ), .op(n9466) );
  nand2_1 U9655 ( .ip1(n12201), .ip2(\cache_data[4][79] ), .op(n9465) );
  nand2_1 U9656 ( .ip1(n12142), .ip2(\cache_data[13][79] ), .op(n9464) );
  nand2_1 U9657 ( .ip1(n9681), .ip2(\cache_data[15][79] ), .op(n9463) );
  nand4_1 U9658 ( .ip1(n9466), .ip2(n9465), .ip3(n9464), .ip4(n9463), .op(
        n9472) );
  nand2_1 U9659 ( .ip1(n9682), .ip2(\cache_data[9][79] ), .op(n9470) );
  nand2_1 U9660 ( .ip1(n9688), .ip2(\cache_data[0][79] ), .op(n9469) );
  nand2_1 U9661 ( .ip1(n9689), .ip2(\cache_data[10][79] ), .op(n9468) );
  nand2_1 U9662 ( .ip1(n9690), .ip2(\cache_data[14][79] ), .op(n9467) );
  nand4_1 U9663 ( .ip1(n9470), .ip2(n9469), .ip3(n9468), .ip4(n9467), .op(
        n9471) );
  nor4_1 U9664 ( .ip1(n9474), .ip2(n9473), .ip3(n9472), .ip4(n9471), .op(
        n11149) );
  nor2_1 U9665 ( .ip1(n11149), .ip2(n10849), .op(n9496) );
  nand2_1 U9666 ( .ip1(n9689), .ip2(\cache_data[10][47] ), .op(n9478) );
  nand2_1 U9667 ( .ip1(n9688), .ip2(\cache_data[0][47] ), .op(n9477) );
  nand2_1 U9668 ( .ip1(n9668), .ip2(\cache_data[8][47] ), .op(n9476) );
  nand2_1 U9669 ( .ip1(n9682), .ip2(\cache_data[9][47] ), .op(n9475) );
  nand4_1 U9670 ( .ip1(n9478), .ip2(n9477), .ip3(n9476), .ip4(n9475), .op(
        n9494) );
  nand2_1 U9671 ( .ip1(n9681), .ip2(\cache_data[15][47] ), .op(n9482) );
  nand2_1 U9672 ( .ip1(n8905), .ip2(\cache_data[6][47] ), .op(n9481) );
  nand2_1 U9673 ( .ip1(n12227), .ip2(\cache_data[12][47] ), .op(n9480) );
  nand2_1 U9674 ( .ip1(n9675), .ip2(\cache_data[5][47] ), .op(n9479) );
  nand4_1 U9675 ( .ip1(n9482), .ip2(n9481), .ip3(n9480), .ip4(n9479), .op(
        n9493) );
  nand2_1 U9676 ( .ip1(n9690), .ip2(\cache_data[14][47] ), .op(n9486) );
  nand2_1 U9677 ( .ip1(n12201), .ip2(\cache_data[4][47] ), .op(n9485) );
  nand2_1 U9678 ( .ip1(n12120), .ip2(\cache_data[1][47] ), .op(n9484) );
  nand2_1 U9679 ( .ip1(n9670), .ip2(\cache_data[7][47] ), .op(n9483) );
  nand4_1 U9680 ( .ip1(n9486), .ip2(n9485), .ip3(n9484), .ip4(n9483), .op(
        n9492) );
  nand2_1 U9681 ( .ip1(n9680), .ip2(\cache_data[3][47] ), .op(n9490) );
  nand2_1 U9682 ( .ip1(n12142), .ip2(\cache_data[13][47] ), .op(n9489) );
  nand2_1 U9683 ( .ip1(n9669), .ip2(\cache_data[11][47] ), .op(n9488) );
  nand2_1 U9684 ( .ip1(n9687), .ip2(\cache_data[2][47] ), .op(n9487) );
  nand4_1 U9685 ( .ip1(n9490), .ip2(n9489), .ip3(n9488), .ip4(n9487), .op(
        n9491) );
  nor4_1 U9686 ( .ip1(n9494), .ip2(n9493), .ip3(n9492), .ip4(n9491), .op(
        n11150) );
  nor2_1 U9687 ( .ip1(n11150), .ip2(n10870), .op(n9495) );
  not_ab_or_c_or_d U9688 ( .ip1(data_wr_mem[15]), .ip2(n10873), .ip3(n9496), 
        .ip4(n9495), .op(n9518) );
  nand2_1 U9689 ( .ip1(n12227), .ip2(\cache_data[12][111] ), .op(n9500) );
  nand2_1 U9690 ( .ip1(n12120), .ip2(\cache_data[1][111] ), .op(n9499) );
  nand2_1 U9691 ( .ip1(n9680), .ip2(\cache_data[3][111] ), .op(n9498) );
  nand2_1 U9692 ( .ip1(n9675), .ip2(\cache_data[5][111] ), .op(n9497) );
  nand4_1 U9693 ( .ip1(n9500), .ip2(n9499), .ip3(n9498), .ip4(n9497), .op(
        n9516) );
  nand2_1 U9694 ( .ip1(n9687), .ip2(\cache_data[2][111] ), .op(n9504) );
  nand2_1 U9695 ( .ip1(n9682), .ip2(\cache_data[9][111] ), .op(n9503) );
  nand2_1 U9696 ( .ip1(n9690), .ip2(\cache_data[14][111] ), .op(n9502) );
  nand2_1 U9697 ( .ip1(n12142), .ip2(\cache_data[13][111] ), .op(n9501) );
  nand4_1 U9698 ( .ip1(n9504), .ip2(n9503), .ip3(n9502), .ip4(n9501), .op(
        n9515) );
  nand2_1 U9699 ( .ip1(n9670), .ip2(\cache_data[7][111] ), .op(n9508) );
  nand2_1 U9700 ( .ip1(n9681), .ip2(\cache_data[15][111] ), .op(n9507) );
  nand2_1 U9701 ( .ip1(n9688), .ip2(\cache_data[0][111] ), .op(n9506) );
  nand2_1 U9702 ( .ip1(n9689), .ip2(\cache_data[10][111] ), .op(n9505) );
  nand4_1 U9703 ( .ip1(n9508), .ip2(n9507), .ip3(n9506), .ip4(n9505), .op(
        n9514) );
  nand2_1 U9704 ( .ip1(n12179), .ip2(\cache_data[6][111] ), .op(n9512) );
  nand2_1 U9705 ( .ip1(n9669), .ip2(\cache_data[11][111] ), .op(n9511) );
  nand2_1 U9706 ( .ip1(n9668), .ip2(\cache_data[8][111] ), .op(n9510) );
  nand2_1 U9707 ( .ip1(n12201), .ip2(\cache_data[4][111] ), .op(n9509) );
  nand4_1 U9708 ( .ip1(n9512), .ip2(n9511), .ip3(n9510), .ip4(n9509), .op(
        n9513) );
  or4_1 U9709 ( .ip1(n9516), .ip2(n9515), .ip3(n9514), .ip4(n9513), .op(n11153) );
  nand2_1 U9710 ( .ip1(n10894), .ip2(n11153), .op(n9517) );
  nand3_1 U9711 ( .ip1(n9519), .ip2(n9518), .ip3(n9517), .op(n7433) );
  nand2_1 U9712 ( .ip1(n9675), .ip2(\cache_data[5][16] ), .op(n9523) );
  nand2_1 U9713 ( .ip1(n9688), .ip2(\cache_data[0][16] ), .op(n9522) );
  nand2_1 U9714 ( .ip1(n9689), .ip2(\cache_data[10][16] ), .op(n9521) );
  nand2_1 U9715 ( .ip1(n12201), .ip2(\cache_data[4][16] ), .op(n9520) );
  nand4_1 U9716 ( .ip1(n9523), .ip2(n9522), .ip3(n9521), .ip4(n9520), .op(
        n9539) );
  nand2_1 U9717 ( .ip1(n9682), .ip2(\cache_data[9][16] ), .op(n9527) );
  nand2_1 U9718 ( .ip1(n12120), .ip2(\cache_data[1][16] ), .op(n9526) );
  nand2_1 U9719 ( .ip1(n9680), .ip2(\cache_data[3][16] ), .op(n9525) );
  nand2_1 U9720 ( .ip1(n12179), .ip2(\cache_data[6][16] ), .op(n9524) );
  nand4_1 U9721 ( .ip1(n9527), .ip2(n9526), .ip3(n9525), .ip4(n9524), .op(
        n9538) );
  nand2_1 U9722 ( .ip1(n9669), .ip2(\cache_data[11][16] ), .op(n9531) );
  nand2_1 U9723 ( .ip1(n9668), .ip2(\cache_data[8][16] ), .op(n9530) );
  nand2_1 U9724 ( .ip1(n12142), .ip2(\cache_data[13][16] ), .op(n9529) );
  nand2_1 U9725 ( .ip1(n9670), .ip2(\cache_data[7][16] ), .op(n9528) );
  nand4_1 U9726 ( .ip1(n9531), .ip2(n9530), .ip3(n9529), .ip4(n9528), .op(
        n9537) );
  nand2_1 U9727 ( .ip1(n9690), .ip2(\cache_data[14][16] ), .op(n9535) );
  nand2_1 U9728 ( .ip1(n9687), .ip2(\cache_data[2][16] ), .op(n9534) );
  nand2_1 U9729 ( .ip1(n9681), .ip2(\cache_data[15][16] ), .op(n9533) );
  nand2_1 U9730 ( .ip1(n12207), .ip2(\cache_data[12][16] ), .op(n9532) );
  nand4_1 U9731 ( .ip1(n9535), .ip2(n9534), .ip3(n9533), .ip4(n9532), .op(
        n9536) );
  or4_1 U9732 ( .ip1(n9539), .ip2(n9538), .ip3(n9537), .ip4(n9536), .op(n11157) );
  nand2_1 U9733 ( .ip1(n10828), .ip2(n11157), .op(n9605) );
  nand2_1 U9734 ( .ip1(n9681), .ip2(\cache_data[15][80] ), .op(n9543) );
  nand2_1 U9735 ( .ip1(n9669), .ip2(\cache_data[11][80] ), .op(n9542) );
  nand2_1 U9736 ( .ip1(n12179), .ip2(\cache_data[6][80] ), .op(n9541) );
  nand2_1 U9737 ( .ip1(n12201), .ip2(\cache_data[4][80] ), .op(n9540) );
  nand4_1 U9738 ( .ip1(n9543), .ip2(n9542), .ip3(n9541), .ip4(n9540), .op(
        n9559) );
  nand2_1 U9739 ( .ip1(n12227), .ip2(\cache_data[12][80] ), .op(n9547) );
  nand2_1 U9740 ( .ip1(n9687), .ip2(\cache_data[2][80] ), .op(n9546) );
  nand2_1 U9741 ( .ip1(n9690), .ip2(\cache_data[14][80] ), .op(n9545) );
  nand2_1 U9742 ( .ip1(n9688), .ip2(\cache_data[0][80] ), .op(n9544) );
  nand4_1 U9743 ( .ip1(n9547), .ip2(n9546), .ip3(n9545), .ip4(n9544), .op(
        n9558) );
  nand2_1 U9744 ( .ip1(n9680), .ip2(\cache_data[3][80] ), .op(n9551) );
  nand2_1 U9745 ( .ip1(n9668), .ip2(\cache_data[8][80] ), .op(n9550) );
  nand2_1 U9746 ( .ip1(n9682), .ip2(\cache_data[9][80] ), .op(n9549) );
  nand2_1 U9747 ( .ip1(n12142), .ip2(\cache_data[13][80] ), .op(n9548) );
  nand4_1 U9748 ( .ip1(n9551), .ip2(n9550), .ip3(n9549), .ip4(n9548), .op(
        n9557) );
  nand2_1 U9749 ( .ip1(n9675), .ip2(\cache_data[5][80] ), .op(n9555) );
  nand2_1 U9750 ( .ip1(n9670), .ip2(\cache_data[7][80] ), .op(n9554) );
  nand2_1 U9751 ( .ip1(n9689), .ip2(\cache_data[10][80] ), .op(n9553) );
  nand2_1 U9752 ( .ip1(n12120), .ip2(\cache_data[1][80] ), .op(n9552) );
  nand4_1 U9753 ( .ip1(n9555), .ip2(n9554), .ip3(n9553), .ip4(n9552), .op(
        n9556) );
  nor4_1 U9754 ( .ip1(n9559), .ip2(n9558), .ip3(n9557), .ip4(n9556), .op(
        n11158) );
  nor2_1 U9755 ( .ip1(n11158), .ip2(n10849), .op(n9582) );
  nand2_1 U9756 ( .ip1(n9689), .ip2(\cache_data[10][48] ), .op(n9564) );
  nand2_1 U9757 ( .ip1(n12142), .ip2(\cache_data[13][48] ), .op(n9563) );
  nand2_1 U9758 ( .ip1(n9560), .ip2(\cache_data[12][48] ), .op(n9562) );
  nand2_1 U9759 ( .ip1(n9682), .ip2(\cache_data[9][48] ), .op(n9561) );
  nand4_1 U9760 ( .ip1(n9564), .ip2(n9563), .ip3(n9562), .ip4(n9561), .op(
        n9580) );
  nand2_1 U9761 ( .ip1(n9669), .ip2(\cache_data[11][48] ), .op(n9568) );
  nand2_1 U9762 ( .ip1(n9690), .ip2(\cache_data[14][48] ), .op(n9567) );
  nand2_1 U9763 ( .ip1(n12120), .ip2(\cache_data[1][48] ), .op(n9566) );
  nand2_1 U9764 ( .ip1(n9668), .ip2(\cache_data[8][48] ), .op(n9565) );
  nand4_1 U9765 ( .ip1(n9568), .ip2(n9567), .ip3(n9566), .ip4(n9565), .op(
        n9579) );
  nand2_1 U9766 ( .ip1(n9670), .ip2(\cache_data[7][48] ), .op(n9572) );
  nand2_1 U9767 ( .ip1(n12201), .ip2(\cache_data[4][48] ), .op(n9571) );
  nand2_1 U9768 ( .ip1(n9687), .ip2(\cache_data[2][48] ), .op(n9570) );
  nand2_1 U9769 ( .ip1(n9681), .ip2(\cache_data[15][48] ), .op(n9569) );
  nand4_1 U9770 ( .ip1(n9572), .ip2(n9571), .ip3(n9570), .ip4(n9569), .op(
        n9578) );
  nand2_1 U9771 ( .ip1(n12179), .ip2(\cache_data[6][48] ), .op(n9576) );
  nand2_1 U9772 ( .ip1(n9680), .ip2(\cache_data[3][48] ), .op(n9575) );
  nand2_1 U9773 ( .ip1(n9688), .ip2(\cache_data[0][48] ), .op(n9574) );
  nand2_1 U9774 ( .ip1(n9675), .ip2(\cache_data[5][48] ), .op(n9573) );
  nand4_1 U9775 ( .ip1(n9576), .ip2(n9575), .ip3(n9574), .ip4(n9573), .op(
        n9577) );
  nor4_1 U9776 ( .ip1(n9580), .ip2(n9579), .ip3(n9578), .ip4(n9577), .op(
        n11159) );
  nor2_1 U9777 ( .ip1(n11159), .ip2(n10870), .op(n9581) );
  not_ab_or_c_or_d U9778 ( .ip1(data_wr_mem[16]), .ip2(n10873), .ip3(n9582), 
        .ip4(n9581), .op(n9604) );
  nand2_1 U9779 ( .ip1(n12120), .ip2(\cache_data[1][112] ), .op(n9586) );
  nand2_1 U9780 ( .ip1(n9681), .ip2(\cache_data[15][112] ), .op(n9585) );
  nand2_1 U9781 ( .ip1(n9675), .ip2(\cache_data[5][112] ), .op(n9584) );
  nand2_1 U9782 ( .ip1(n9687), .ip2(\cache_data[2][112] ), .op(n9583) );
  nand4_1 U9783 ( .ip1(n9586), .ip2(n9585), .ip3(n9584), .ip4(n9583), .op(
        n9602) );
  nand2_1 U9784 ( .ip1(n9682), .ip2(\cache_data[9][112] ), .op(n9590) );
  nand2_1 U9785 ( .ip1(n9688), .ip2(\cache_data[0][112] ), .op(n9589) );
  nand2_1 U9786 ( .ip1(n12142), .ip2(\cache_data[13][112] ), .op(n9588) );
  nand2_1 U9787 ( .ip1(n9689), .ip2(\cache_data[10][112] ), .op(n9587) );
  nand4_1 U9788 ( .ip1(n9590), .ip2(n9589), .ip3(n9588), .ip4(n9587), .op(
        n9601) );
  nand2_1 U9789 ( .ip1(n12227), .ip2(\cache_data[12][112] ), .op(n9594) );
  nand2_1 U9790 ( .ip1(n9670), .ip2(\cache_data[7][112] ), .op(n9593) );
  nand2_1 U9791 ( .ip1(n9690), .ip2(\cache_data[14][112] ), .op(n9592) );
  nand2_1 U9792 ( .ip1(n12179), .ip2(\cache_data[6][112] ), .op(n9591) );
  nand4_1 U9793 ( .ip1(n9594), .ip2(n9593), .ip3(n9592), .ip4(n9591), .op(
        n9600) );
  nand2_1 U9794 ( .ip1(n9668), .ip2(\cache_data[8][112] ), .op(n9598) );
  nand2_1 U9795 ( .ip1(n9669), .ip2(\cache_data[11][112] ), .op(n9597) );
  nand2_1 U9796 ( .ip1(n12201), .ip2(\cache_data[4][112] ), .op(n9596) );
  nand2_1 U9797 ( .ip1(n9680), .ip2(\cache_data[3][112] ), .op(n9595) );
  nand4_1 U9798 ( .ip1(n9598), .ip2(n9597), .ip3(n9596), .ip4(n9595), .op(
        n9599) );
  or4_1 U9799 ( .ip1(n9602), .ip2(n9601), .ip3(n9600), .ip4(n9599), .op(n11162) );
  nand2_1 U9800 ( .ip1(n10894), .ip2(n11162), .op(n9603) );
  nand3_1 U9801 ( .ip1(n9605), .ip2(n9604), .ip3(n9603), .op(n7432) );
  nand2_1 U9802 ( .ip1(data_wr_mem[17]), .ip2(n10873), .op(n9701) );
  nand2_1 U9803 ( .ip1(n12227), .ip2(\cache_data[12][113] ), .op(n9609) );
  nand2_1 U9804 ( .ip1(n9680), .ip2(\cache_data[3][113] ), .op(n9608) );
  nand2_1 U9805 ( .ip1(n12120), .ip2(\cache_data[1][113] ), .op(n9607) );
  nand2_1 U9806 ( .ip1(n9681), .ip2(\cache_data[15][113] ), .op(n9606) );
  nand4_1 U9807 ( .ip1(n9609), .ip2(n9608), .ip3(n9607), .ip4(n9606), .op(
        n9625) );
  nand2_1 U9808 ( .ip1(n9690), .ip2(\cache_data[14][113] ), .op(n9613) );
  nand2_1 U9809 ( .ip1(n9669), .ip2(\cache_data[11][113] ), .op(n9612) );
  nand2_1 U9810 ( .ip1(n9687), .ip2(\cache_data[2][113] ), .op(n9611) );
  nand2_1 U9811 ( .ip1(n12201), .ip2(\cache_data[4][113] ), .op(n9610) );
  nand4_1 U9812 ( .ip1(n9613), .ip2(n9612), .ip3(n9611), .ip4(n9610), .op(
        n9624) );
  nand2_1 U9813 ( .ip1(n9668), .ip2(\cache_data[8][113] ), .op(n9617) );
  nand2_1 U9814 ( .ip1(n9675), .ip2(\cache_data[5][113] ), .op(n9616) );
  nand2_1 U9815 ( .ip1(n9689), .ip2(\cache_data[10][113] ), .op(n9615) );
  nand2_1 U9816 ( .ip1(n9682), .ip2(\cache_data[9][113] ), .op(n9614) );
  nand4_1 U9817 ( .ip1(n9617), .ip2(n9616), .ip3(n9615), .ip4(n9614), .op(
        n9623) );
  nand2_1 U9818 ( .ip1(n9670), .ip2(\cache_data[7][113] ), .op(n9621) );
  nand2_1 U9819 ( .ip1(n12142), .ip2(\cache_data[13][113] ), .op(n9620) );
  nand2_1 U9820 ( .ip1(n12179), .ip2(\cache_data[6][113] ), .op(n9619) );
  nand2_1 U9821 ( .ip1(n9688), .ip2(\cache_data[0][113] ), .op(n9618) );
  nand4_1 U9822 ( .ip1(n9621), .ip2(n9620), .ip3(n9619), .ip4(n9618), .op(
        n9622) );
  or4_1 U9823 ( .ip1(n9625), .ip2(n9624), .ip3(n9623), .ip4(n9622), .op(n11166) );
  nand2_1 U9824 ( .ip1(n9682), .ip2(\cache_data[9][81] ), .op(n9629) );
  nand2_1 U9825 ( .ip1(n9681), .ip2(\cache_data[15][81] ), .op(n9628) );
  nand2_1 U9826 ( .ip1(n12227), .ip2(\cache_data[12][81] ), .op(n9627) );
  nand2_1 U9827 ( .ip1(n9680), .ip2(\cache_data[3][81] ), .op(n9626) );
  nand4_1 U9828 ( .ip1(n9629), .ip2(n9628), .ip3(n9627), .ip4(n9626), .op(
        n9645) );
  nand2_1 U9829 ( .ip1(n9669), .ip2(\cache_data[11][81] ), .op(n9633) );
  nand2_1 U9830 ( .ip1(n12179), .ip2(\cache_data[6][81] ), .op(n9632) );
  nand2_1 U9831 ( .ip1(n9690), .ip2(\cache_data[14][81] ), .op(n9631) );
  nand2_1 U9832 ( .ip1(n12242), .ip2(\cache_data[13][81] ), .op(n9630) );
  nand4_1 U9833 ( .ip1(n9633), .ip2(n9632), .ip3(n9631), .ip4(n9630), .op(
        n9644) );
  nand2_1 U9834 ( .ip1(n9687), .ip2(\cache_data[2][81] ), .op(n9637) );
  nand2_1 U9835 ( .ip1(n9675), .ip2(\cache_data[5][81] ), .op(n9636) );
  nand2_1 U9836 ( .ip1(n9689), .ip2(\cache_data[10][81] ), .op(n9635) );
  nand2_1 U9837 ( .ip1(n9688), .ip2(\cache_data[0][81] ), .op(n9634) );
  nand4_1 U9838 ( .ip1(n9637), .ip2(n9636), .ip3(n9635), .ip4(n9634), .op(
        n9643) );
  nand2_1 U9839 ( .ip1(n9670), .ip2(\cache_data[7][81] ), .op(n9641) );
  nand2_1 U9840 ( .ip1(n8906), .ip2(\cache_data[4][81] ), .op(n9640) );
  nand2_1 U9841 ( .ip1(n9668), .ip2(\cache_data[8][81] ), .op(n9639) );
  nand2_1 U9842 ( .ip1(n12120), .ip2(\cache_data[1][81] ), .op(n9638) );
  nand4_1 U9843 ( .ip1(n9641), .ip2(n9640), .ip3(n9639), .ip4(n9638), .op(
        n9642) );
  nor4_1 U9844 ( .ip1(n9645), .ip2(n9644), .ip3(n9643), .ip4(n9642), .op(
        n11168) );
  nor2_1 U9845 ( .ip1(n11168), .ip2(n10849), .op(n9667) );
  nand2_1 U9846 ( .ip1(n9670), .ip2(\cache_data[7][49] ), .op(n9649) );
  nand2_1 U9847 ( .ip1(n12142), .ip2(\cache_data[13][49] ), .op(n9648) );
  nand2_1 U9848 ( .ip1(n9669), .ip2(\cache_data[11][49] ), .op(n9647) );
  nand2_1 U9849 ( .ip1(n9690), .ip2(\cache_data[14][49] ), .op(n9646) );
  nand4_1 U9850 ( .ip1(n9649), .ip2(n9648), .ip3(n9647), .ip4(n9646), .op(
        n9665) );
  nand2_1 U9851 ( .ip1(n12243), .ip2(\cache_data[4][49] ), .op(n9653) );
  nand2_1 U9852 ( .ip1(n9682), .ip2(\cache_data[9][49] ), .op(n9652) );
  nand2_1 U9853 ( .ip1(n12227), .ip2(\cache_data[12][49] ), .op(n9651) );
  nand2_1 U9854 ( .ip1(n9675), .ip2(\cache_data[5][49] ), .op(n9650) );
  nand4_1 U9855 ( .ip1(n9653), .ip2(n9652), .ip3(n9651), .ip4(n9650), .op(
        n9664) );
  nand2_1 U9856 ( .ip1(n9668), .ip2(\cache_data[8][49] ), .op(n9657) );
  nand2_1 U9857 ( .ip1(n9687), .ip2(\cache_data[2][49] ), .op(n9656) );
  nand2_1 U9858 ( .ip1(n9688), .ip2(\cache_data[0][49] ), .op(n9655) );
  nand2_1 U9859 ( .ip1(n12120), .ip2(\cache_data[1][49] ), .op(n9654) );
  nand4_1 U9860 ( .ip1(n9657), .ip2(n9656), .ip3(n9655), .ip4(n9654), .op(
        n9663) );
  nand2_1 U9861 ( .ip1(n9689), .ip2(\cache_data[10][49] ), .op(n9661) );
  nand2_1 U9862 ( .ip1(n9681), .ip2(\cache_data[15][49] ), .op(n9660) );
  nand2_1 U9863 ( .ip1(n12179), .ip2(\cache_data[6][49] ), .op(n9659) );
  nand2_1 U9864 ( .ip1(n9680), .ip2(\cache_data[3][49] ), .op(n9658) );
  nand4_1 U9865 ( .ip1(n9661), .ip2(n9660), .ip3(n9659), .ip4(n9658), .op(
        n9662) );
  nor4_1 U9866 ( .ip1(n9665), .ip2(n9664), .ip3(n9663), .ip4(n9662), .op(
        n11167) );
  nor2_1 U9867 ( .ip1(n11167), .ip2(n10870), .op(n9666) );
  not_ab_or_c_or_d U9868 ( .ip1(n10894), .ip2(n11166), .ip3(n9667), .ip4(n9666), .op(n9700) );
  nand2_1 U9869 ( .ip1(n9668), .ip2(\cache_data[8][17] ), .op(n9674) );
  nand2_1 U9870 ( .ip1(n9669), .ip2(\cache_data[11][17] ), .op(n9673) );
  nand2_1 U9871 ( .ip1(n9670), .ip2(\cache_data[7][17] ), .op(n9672) );
  nand2_1 U9872 ( .ip1(n12179), .ip2(\cache_data[6][17] ), .op(n9671) );
  nand4_1 U9873 ( .ip1(n9674), .ip2(n9673), .ip3(n9672), .ip4(n9671), .op(
        n9698) );
  nand2_1 U9874 ( .ip1(n12142), .ip2(\cache_data[13][17] ), .op(n9679) );
  nand2_1 U9875 ( .ip1(n12207), .ip2(\cache_data[12][17] ), .op(n9678) );
  nand2_1 U9876 ( .ip1(n12120), .ip2(\cache_data[1][17] ), .op(n9677) );
  nand2_1 U9877 ( .ip1(n9675), .ip2(\cache_data[5][17] ), .op(n9676) );
  nand4_1 U9878 ( .ip1(n9679), .ip2(n9678), .ip3(n9677), .ip4(n9676), .op(
        n9697) );
  nand2_1 U9879 ( .ip1(n9680), .ip2(\cache_data[3][17] ), .op(n9686) );
  nand2_1 U9880 ( .ip1(n9681), .ip2(\cache_data[15][17] ), .op(n9685) );
  nand2_1 U9881 ( .ip1(n12201), .ip2(\cache_data[4][17] ), .op(n9684) );
  nand2_1 U9882 ( .ip1(n9682), .ip2(\cache_data[9][17] ), .op(n9683) );
  nand4_1 U9883 ( .ip1(n9686), .ip2(n9685), .ip3(n9684), .ip4(n9683), .op(
        n9696) );
  nand2_1 U9884 ( .ip1(n9687), .ip2(\cache_data[2][17] ), .op(n9694) );
  nand2_1 U9885 ( .ip1(n9688), .ip2(\cache_data[0][17] ), .op(n9693) );
  nand2_1 U9886 ( .ip1(n9689), .ip2(\cache_data[10][17] ), .op(n9692) );
  nand2_1 U9887 ( .ip1(n9690), .ip2(\cache_data[14][17] ), .op(n9691) );
  nand4_1 U9888 ( .ip1(n9694), .ip2(n9693), .ip3(n9692), .ip4(n9691), .op(
        n9695) );
  or4_1 U9889 ( .ip1(n9698), .ip2(n9697), .ip3(n9696), .ip4(n9695), .op(n11171) );
  nand2_1 U9890 ( .ip1(n10828), .ip2(n11171), .op(n9699) );
  nand3_1 U9891 ( .ip1(n9701), .ip2(n9700), .ip3(n9699), .op(n7431) );
  nand2_1 U9892 ( .ip1(data_wr_mem[18]), .ip2(n10873), .op(n9786) );
  nand2_1 U9893 ( .ip1(n12243), .ip2(\cache_data[4][114] ), .op(n9705) );
  nand2_1 U9894 ( .ip1(n12165), .ip2(\cache_data[13][114] ), .op(n9704) );
  nand2_1 U9895 ( .ip1(n12191), .ip2(\cache_data[8][114] ), .op(n9703) );
  nand2_1 U9896 ( .ip1(n12179), .ip2(\cache_data[6][114] ), .op(n9702) );
  nand4_1 U9897 ( .ip1(n9705), .ip2(n9704), .ip3(n9703), .ip4(n9702), .op(
        n9721) );
  nand2_1 U9898 ( .ip1(n12202), .ip2(\cache_data[7][114] ), .op(n9709) );
  nand2_1 U9899 ( .ip1(n12233), .ip2(\cache_data[0][114] ), .op(n9708) );
  nand2_1 U9900 ( .ip1(n12219), .ip2(\cache_data[3][114] ), .op(n9707) );
  nand2_1 U9901 ( .ip1(n11927), .ip2(\cache_data[11][114] ), .op(n9706) );
  nand4_1 U9902 ( .ip1(n9709), .ip2(n9708), .ip3(n9707), .ip4(n9706), .op(
        n9720) );
  nand2_1 U9903 ( .ip1(n12228), .ip2(\cache_data[2][114] ), .op(n9713) );
  nand2_1 U9904 ( .ip1(n12240), .ip2(\cache_data[5][114] ), .op(n9712) );
  nand2_1 U9905 ( .ip1(n12221), .ip2(\cache_data[15][114] ), .op(n9711) );
  nand2_1 U9906 ( .ip1(n12227), .ip2(\cache_data[12][114] ), .op(n9710) );
  nand4_1 U9907 ( .ip1(n9713), .ip2(n9712), .ip3(n9711), .ip4(n9710), .op(
        n9719) );
  nand2_1 U9908 ( .ip1(n12220), .ip2(\cache_data[14][114] ), .op(n9717) );
  nand2_1 U9909 ( .ip1(n12235), .ip2(\cache_data[10][114] ), .op(n9716) );
  nand2_1 U9910 ( .ip1(n8894), .ip2(\cache_data[1][114] ), .op(n9715) );
  nand2_1 U9911 ( .ip1(n12241), .ip2(\cache_data[9][114] ), .op(n9714) );
  nand4_1 U9912 ( .ip1(n9717), .ip2(n9716), .ip3(n9715), .ip4(n9714), .op(
        n9718) );
  or4_1 U9913 ( .ip1(n9721), .ip2(n9720), .ip3(n9719), .ip4(n9718), .op(n11180) );
  nand2_1 U9914 ( .ip1(n12241), .ip2(\cache_data[9][82] ), .op(n9725) );
  nand2_1 U9915 ( .ip1(n12220), .ip2(\cache_data[14][82] ), .op(n9724) );
  nand2_1 U9916 ( .ip1(n12191), .ip2(\cache_data[8][82] ), .op(n9723) );
  nand2_1 U9917 ( .ip1(n12233), .ip2(\cache_data[0][82] ), .op(n9722) );
  nand4_1 U9918 ( .ip1(n9725), .ip2(n9724), .ip3(n9723), .ip4(n9722), .op(
        n9741) );
  nand2_1 U9919 ( .ip1(n12235), .ip2(\cache_data[10][82] ), .op(n9729) );
  nand2_1 U9920 ( .ip1(n8894), .ip2(\cache_data[1][82] ), .op(n9728) );
  nand2_1 U9921 ( .ip1(n11927), .ip2(\cache_data[11][82] ), .op(n9727) );
  nand2_1 U9922 ( .ip1(n12228), .ip2(\cache_data[2][82] ), .op(n9726) );
  nand4_1 U9923 ( .ip1(n9729), .ip2(n9728), .ip3(n9727), .ip4(n9726), .op(
        n9740) );
  nand2_1 U9924 ( .ip1(n12221), .ip2(\cache_data[15][82] ), .op(n9733) );
  nand2_1 U9925 ( .ip1(n12243), .ip2(\cache_data[4][82] ), .op(n9732) );
  nand2_1 U9926 ( .ip1(n12165), .ip2(\cache_data[13][82] ), .op(n9731) );
  nand2_1 U9927 ( .ip1(n12179), .ip2(\cache_data[6][82] ), .op(n9730) );
  nand4_1 U9928 ( .ip1(n9733), .ip2(n9732), .ip3(n9731), .ip4(n9730), .op(
        n9739) );
  nand2_1 U9929 ( .ip1(n12227), .ip2(\cache_data[12][82] ), .op(n9737) );
  nand2_1 U9930 ( .ip1(n12219), .ip2(\cache_data[3][82] ), .op(n9736) );
  nand2_1 U9931 ( .ip1(n12202), .ip2(\cache_data[7][82] ), .op(n9735) );
  nand2_1 U9932 ( .ip1(n12240), .ip2(\cache_data[5][82] ), .op(n9734) );
  nand4_1 U9933 ( .ip1(n9737), .ip2(n9736), .ip3(n9735), .ip4(n9734), .op(
        n9738) );
  nor4_1 U9934 ( .ip1(n9741), .ip2(n9740), .ip3(n9739), .ip4(n9738), .op(
        n11177) );
  nor2_1 U9935 ( .ip1(n11177), .ip2(n10849), .op(n9763) );
  nand2_1 U9936 ( .ip1(n12179), .ip2(\cache_data[6][50] ), .op(n9745) );
  nand2_1 U9937 ( .ip1(n12235), .ip2(\cache_data[10][50] ), .op(n9744) );
  nand2_1 U9938 ( .ip1(n12243), .ip2(\cache_data[4][50] ), .op(n9743) );
  nand2_1 U9939 ( .ip1(n12202), .ip2(\cache_data[7][50] ), .op(n9742) );
  nand4_1 U9940 ( .ip1(n9745), .ip2(n9744), .ip3(n9743), .ip4(n9742), .op(
        n9761) );
  nand2_1 U9941 ( .ip1(n12233), .ip2(\cache_data[0][50] ), .op(n9749) );
  nand2_1 U9942 ( .ip1(n12240), .ip2(\cache_data[5][50] ), .op(n9748) );
  nand2_1 U9943 ( .ip1(n11971), .ip2(\cache_data[14][50] ), .op(n9747) );
  nand2_1 U9944 ( .ip1(n12219), .ip2(\cache_data[3][50] ), .op(n9746) );
  nand4_1 U9945 ( .ip1(n9749), .ip2(n9748), .ip3(n9747), .ip4(n9746), .op(
        n9760) );
  nand2_1 U9946 ( .ip1(n12221), .ip2(\cache_data[15][50] ), .op(n9753) );
  nand2_1 U9947 ( .ip1(n12227), .ip2(\cache_data[12][50] ), .op(n9752) );
  nand2_1 U9948 ( .ip1(n11927), .ip2(\cache_data[11][50] ), .op(n9751) );
  nand2_1 U9949 ( .ip1(n12191), .ip2(\cache_data[8][50] ), .op(n9750) );
  nand4_1 U9950 ( .ip1(n9753), .ip2(n9752), .ip3(n9751), .ip4(n9750), .op(
        n9759) );
  nand2_1 U9951 ( .ip1(n12165), .ip2(\cache_data[13][50] ), .op(n9757) );
  nand2_1 U9952 ( .ip1(n12241), .ip2(\cache_data[9][50] ), .op(n9756) );
  nand2_1 U9953 ( .ip1(n8894), .ip2(\cache_data[1][50] ), .op(n9755) );
  nand2_1 U9954 ( .ip1(n12228), .ip2(\cache_data[2][50] ), .op(n9754) );
  nand4_1 U9955 ( .ip1(n9757), .ip2(n9756), .ip3(n9755), .ip4(n9754), .op(
        n9758) );
  nor4_1 U9956 ( .ip1(n9761), .ip2(n9760), .ip3(n9759), .ip4(n9758), .op(
        n11176) );
  nor2_1 U9957 ( .ip1(n11176), .ip2(n10870), .op(n9762) );
  not_ab_or_c_or_d U9958 ( .ip1(n10894), .ip2(n11180), .ip3(n9763), .ip4(n9762), .op(n9785) );
  nand2_1 U9959 ( .ip1(n12221), .ip2(\cache_data[15][18] ), .op(n9767) );
  nand2_1 U9960 ( .ip1(n11943), .ip2(\cache_data[1][18] ), .op(n9766) );
  nand2_1 U9961 ( .ip1(n12201), .ip2(\cache_data[4][18] ), .op(n9765) );
  nand2_1 U9962 ( .ip1(n12235), .ip2(\cache_data[10][18] ), .op(n9764) );
  nand4_1 U9963 ( .ip1(n9767), .ip2(n9766), .ip3(n9765), .ip4(n9764), .op(
        n9783) );
  nand2_1 U9964 ( .ip1(n12126), .ip2(\cache_data[9][18] ), .op(n9771) );
  nand2_1 U9965 ( .ip1(n12226), .ip2(\cache_data[7][18] ), .op(n9770) );
  nand2_1 U9966 ( .ip1(n12228), .ip2(\cache_data[2][18] ), .op(n9769) );
  nand2_1 U9967 ( .ip1(n12233), .ip2(\cache_data[0][18] ), .op(n9768) );
  nand4_1 U9968 ( .ip1(n9771), .ip2(n9770), .ip3(n9769), .ip4(n9768), .op(
        n9782) );
  nand2_1 U9969 ( .ip1(n12179), .ip2(\cache_data[6][18] ), .op(n9775) );
  nand2_1 U9970 ( .ip1(n12219), .ip2(\cache_data[3][18] ), .op(n9774) );
  nand2_1 U9971 ( .ip1(n12240), .ip2(\cache_data[5][18] ), .op(n9773) );
  nand2_1 U9972 ( .ip1(n12142), .ip2(\cache_data[13][18] ), .op(n9772) );
  nand4_1 U9973 ( .ip1(n9775), .ip2(n9774), .ip3(n9773), .ip4(n9772), .op(
        n9781) );
  nand2_1 U9974 ( .ip1(n12220), .ip2(\cache_data[14][18] ), .op(n9779) );
  nand2_1 U9975 ( .ip1(n12121), .ip2(\cache_data[8][18] ), .op(n9778) );
  nand2_1 U9976 ( .ip1(n12207), .ip2(\cache_data[12][18] ), .op(n9777) );
  nand2_1 U9977 ( .ip1(n12096), .ip2(\cache_data[11][18] ), .op(n9776) );
  nand4_1 U9978 ( .ip1(n9779), .ip2(n9778), .ip3(n9777), .ip4(n9776), .op(
        n9780) );
  or4_1 U9979 ( .ip1(n9783), .ip2(n9782), .ip3(n9781), .ip4(n9780), .op(n11175) );
  nand2_1 U9980 ( .ip1(n10828), .ip2(n11175), .op(n9784) );
  nand3_1 U9981 ( .ip1(n9786), .ip2(n9785), .ip3(n9784), .op(n7430) );
  nand2_1 U9982 ( .ip1(n12179), .ip2(\cache_data[6][19] ), .op(n9790) );
  nand2_1 U9983 ( .ip1(n12201), .ip2(\cache_data[4][19] ), .op(n9789) );
  nand2_1 U9984 ( .ip1(n12219), .ip2(\cache_data[3][19] ), .op(n9788) );
  nand2_1 U9985 ( .ip1(n12142), .ip2(\cache_data[13][19] ), .op(n9787) );
  nand4_1 U9986 ( .ip1(n9790), .ip2(n9789), .ip3(n9788), .ip4(n9787), .op(
        n9806) );
  nand2_1 U9987 ( .ip1(n12121), .ip2(\cache_data[8][19] ), .op(n9794) );
  nand2_1 U9988 ( .ip1(n12233), .ip2(\cache_data[0][19] ), .op(n9793) );
  nand2_1 U9989 ( .ip1(n12240), .ip2(\cache_data[5][19] ), .op(n9792) );
  nand2_1 U9990 ( .ip1(n12220), .ip2(\cache_data[14][19] ), .op(n9791) );
  nand4_1 U9991 ( .ip1(n9794), .ip2(n9793), .ip3(n9792), .ip4(n9791), .op(
        n9805) );
  nand2_1 U9992 ( .ip1(n11943), .ip2(\cache_data[1][19] ), .op(n9798) );
  nand2_1 U9993 ( .ip1(n12228), .ip2(\cache_data[2][19] ), .op(n9797) );
  nand2_1 U9994 ( .ip1(n12235), .ip2(\cache_data[10][19] ), .op(n9796) );
  nand2_1 U9995 ( .ip1(n12096), .ip2(\cache_data[11][19] ), .op(n9795) );
  nand4_1 U9996 ( .ip1(n9798), .ip2(n9797), .ip3(n9796), .ip4(n9795), .op(
        n9804) );
  nand2_1 U9997 ( .ip1(n12226), .ip2(\cache_data[7][19] ), .op(n9802) );
  nand2_1 U9998 ( .ip1(n12126), .ip2(\cache_data[9][19] ), .op(n9801) );
  nand2_1 U9999 ( .ip1(n12221), .ip2(\cache_data[15][19] ), .op(n9800) );
  nand2_1 U10000 ( .ip1(n12207), .ip2(\cache_data[12][19] ), .op(n9799) );
  nand4_1 U10001 ( .ip1(n9802), .ip2(n9801), .ip3(n9800), .ip4(n9799), .op(
        n9803) );
  or4_1 U10002 ( .ip1(n9806), .ip2(n9805), .ip3(n9804), .ip4(n9803), .op(
        n11184) );
  nand2_1 U10003 ( .ip1(n10828), .ip2(n11184), .op(n9871) );
  nand2_1 U10004 ( .ip1(n12179), .ip2(\cache_data[6][83] ), .op(n9810) );
  nand2_1 U10005 ( .ip1(n12227), .ip2(\cache_data[12][83] ), .op(n9809) );
  nand2_1 U10006 ( .ip1(n12219), .ip2(\cache_data[3][83] ), .op(n9808) );
  nand2_1 U10007 ( .ip1(n12235), .ip2(\cache_data[10][83] ), .op(n9807) );
  nand4_1 U10008 ( .ip1(n9810), .ip2(n9809), .ip3(n9808), .ip4(n9807), .op(
        n9826) );
  nand2_1 U10009 ( .ip1(n12165), .ip2(\cache_data[13][83] ), .op(n9814) );
  nand2_1 U10010 ( .ip1(n8894), .ip2(\cache_data[1][83] ), .op(n9813) );
  nand2_1 U10011 ( .ip1(n12243), .ip2(\cache_data[4][83] ), .op(n9812) );
  nand2_1 U10012 ( .ip1(n11927), .ip2(\cache_data[11][83] ), .op(n9811) );
  nand4_1 U10013 ( .ip1(n9814), .ip2(n9813), .ip3(n9812), .ip4(n9811), .op(
        n9825) );
  nand2_1 U10014 ( .ip1(n12221), .ip2(\cache_data[15][83] ), .op(n9818) );
  nand2_1 U10015 ( .ip1(n12233), .ip2(\cache_data[0][83] ), .op(n9817) );
  nand2_1 U10016 ( .ip1(n12202), .ip2(\cache_data[7][83] ), .op(n9816) );
  nand2_1 U10017 ( .ip1(n12240), .ip2(\cache_data[5][83] ), .op(n9815) );
  nand4_1 U10018 ( .ip1(n9818), .ip2(n9817), .ip3(n9816), .ip4(n9815), .op(
        n9824) );
  nand2_1 U10019 ( .ip1(n12241), .ip2(\cache_data[9][83] ), .op(n9822) );
  nand2_1 U10020 ( .ip1(n12191), .ip2(\cache_data[8][83] ), .op(n9821) );
  nand2_1 U10021 ( .ip1(n12220), .ip2(\cache_data[14][83] ), .op(n9820) );
  nand2_1 U10022 ( .ip1(n12228), .ip2(\cache_data[2][83] ), .op(n9819) );
  nand4_1 U10023 ( .ip1(n9822), .ip2(n9821), .ip3(n9820), .ip4(n9819), .op(
        n9823) );
  nor4_1 U10024 ( .ip1(n9826), .ip2(n9825), .ip3(n9824), .ip4(n9823), .op(
        n11185) );
  nor2_1 U10025 ( .ip1(n11185), .ip2(n10849), .op(n9848) );
  nand2_1 U10026 ( .ip1(n12243), .ip2(\cache_data[4][51] ), .op(n9830) );
  nand2_1 U10027 ( .ip1(n12202), .ip2(\cache_data[7][51] ), .op(n9829) );
  nand2_1 U10028 ( .ip1(n12241), .ip2(\cache_data[9][51] ), .op(n9828) );
  nand2_1 U10029 ( .ip1(n12219), .ip2(\cache_data[3][51] ), .op(n9827) );
  nand4_1 U10030 ( .ip1(n9830), .ip2(n9829), .ip3(n9828), .ip4(n9827), .op(
        n9846) );
  nand2_1 U10031 ( .ip1(n12179), .ip2(\cache_data[6][51] ), .op(n9834) );
  nand2_1 U10032 ( .ip1(n11927), .ip2(\cache_data[11][51] ), .op(n9833) );
  nand2_1 U10033 ( .ip1(n12191), .ip2(\cache_data[8][51] ), .op(n9832) );
  nand2_1 U10034 ( .ip1(n12235), .ip2(\cache_data[10][51] ), .op(n9831) );
  nand4_1 U10035 ( .ip1(n9834), .ip2(n9833), .ip3(n9832), .ip4(n9831), .op(
        n9845) );
  nand2_1 U10036 ( .ip1(n12233), .ip2(\cache_data[0][51] ), .op(n9838) );
  nand2_1 U10037 ( .ip1(n12240), .ip2(\cache_data[5][51] ), .op(n9837) );
  nand2_1 U10038 ( .ip1(n12227), .ip2(\cache_data[12][51] ), .op(n9836) );
  nand2_1 U10039 ( .ip1(n12221), .ip2(\cache_data[15][51] ), .op(n9835) );
  nand4_1 U10040 ( .ip1(n9838), .ip2(n9837), .ip3(n9836), .ip4(n9835), .op(
        n9844) );
  nand2_1 U10041 ( .ip1(n12220), .ip2(\cache_data[14][51] ), .op(n9842) );
  nand2_1 U10042 ( .ip1(n8894), .ip2(\cache_data[1][51] ), .op(n9841) );
  nand2_1 U10043 ( .ip1(n12165), .ip2(\cache_data[13][51] ), .op(n9840) );
  nand2_1 U10044 ( .ip1(n12228), .ip2(\cache_data[2][51] ), .op(n9839) );
  nand4_1 U10045 ( .ip1(n9842), .ip2(n9841), .ip3(n9840), .ip4(n9839), .op(
        n9843) );
  nor4_1 U10046 ( .ip1(n9846), .ip2(n9845), .ip3(n9844), .ip4(n9843), .op(
        n11186) );
  nor2_1 U10047 ( .ip1(n11186), .ip2(n10870), .op(n9847) );
  not_ab_or_c_or_d U10048 ( .ip1(data_wr_mem[19]), .ip2(n10873), .ip3(n9848), 
        .ip4(n9847), .op(n9870) );
  nand2_1 U10049 ( .ip1(n12121), .ip2(\cache_data[8][115] ), .op(n9852) );
  nand2_1 U10050 ( .ip1(n12221), .ip2(\cache_data[15][115] ), .op(n9851) );
  nand2_1 U10051 ( .ip1(n12235), .ip2(\cache_data[10][115] ), .op(n9850) );
  nand2_1 U10052 ( .ip1(n12219), .ip2(\cache_data[3][115] ), .op(n9849) );
  nand4_1 U10053 ( .ip1(n9852), .ip2(n9851), .ip3(n9850), .ip4(n9849), .op(
        n9868) );
  nand2_1 U10054 ( .ip1(n12240), .ip2(\cache_data[5][115] ), .op(n9856) );
  nand2_1 U10055 ( .ip1(n12142), .ip2(\cache_data[13][115] ), .op(n9855) );
  nand2_1 U10056 ( .ip1(n12226), .ip2(\cache_data[7][115] ), .op(n9854) );
  nand2_1 U10057 ( .ip1(n12207), .ip2(\cache_data[12][115] ), .op(n9853) );
  nand4_1 U10058 ( .ip1(n9856), .ip2(n9855), .ip3(n9854), .ip4(n9853), .op(
        n9867) );
  nand2_1 U10059 ( .ip1(n12201), .ip2(\cache_data[4][115] ), .op(n9860) );
  nand2_1 U10060 ( .ip1(n11979), .ip2(\cache_data[1][115] ), .op(n9859) );
  nand2_1 U10061 ( .ip1(n12228), .ip2(\cache_data[2][115] ), .op(n9858) );
  nand2_1 U10062 ( .ip1(n12220), .ip2(\cache_data[14][115] ), .op(n9857) );
  nand4_1 U10063 ( .ip1(n9860), .ip2(n9859), .ip3(n9858), .ip4(n9857), .op(
        n9866) );
  nand2_1 U10064 ( .ip1(n12179), .ip2(\cache_data[6][115] ), .op(n9864) );
  nand2_1 U10065 ( .ip1(n12233), .ip2(\cache_data[0][115] ), .op(n9863) );
  nand2_1 U10066 ( .ip1(n12096), .ip2(\cache_data[11][115] ), .op(n9862) );
  nand2_1 U10067 ( .ip1(n12126), .ip2(\cache_data[9][115] ), .op(n9861) );
  nand4_1 U10068 ( .ip1(n9864), .ip2(n9863), .ip3(n9862), .ip4(n9861), .op(
        n9865) );
  or4_1 U10069 ( .ip1(n9868), .ip2(n9867), .ip3(n9866), .ip4(n9865), .op(
        n11189) );
  nand2_1 U10070 ( .ip1(n10894), .ip2(n11189), .op(n9869) );
  nand3_1 U10071 ( .ip1(n9871), .ip2(n9870), .ip3(n9869), .op(n7429) );
  nand2_1 U10072 ( .ip1(n12235), .ip2(\cache_data[10][20] ), .op(n9875) );
  nand2_1 U10073 ( .ip1(n12220), .ip2(\cache_data[14][20] ), .op(n9874) );
  nand2_1 U10074 ( .ip1(n12126), .ip2(\cache_data[9][20] ), .op(n9873) );
  nand2_1 U10075 ( .ip1(n12179), .ip2(\cache_data[6][20] ), .op(n9872) );
  nand4_1 U10076 ( .ip1(n9875), .ip2(n9874), .ip3(n9873), .ip4(n9872), .op(
        n9891) );
  nand2_1 U10077 ( .ip1(n12121), .ip2(\cache_data[8][20] ), .op(n9879) );
  nand2_1 U10078 ( .ip1(n11979), .ip2(\cache_data[1][20] ), .op(n9878) );
  nand2_1 U10079 ( .ip1(n12228), .ip2(\cache_data[2][20] ), .op(n9877) );
  nand2_1 U10080 ( .ip1(n12142), .ip2(\cache_data[13][20] ), .op(n9876) );
  nand4_1 U10081 ( .ip1(n9879), .ip2(n9878), .ip3(n9877), .ip4(n9876), .op(
        n9890) );
  nand2_1 U10082 ( .ip1(n12207), .ip2(\cache_data[12][20] ), .op(n9883) );
  nand2_1 U10083 ( .ip1(n12219), .ip2(\cache_data[3][20] ), .op(n9882) );
  nand2_1 U10084 ( .ip1(n12233), .ip2(\cache_data[0][20] ), .op(n9881) );
  nand2_1 U10085 ( .ip1(n12240), .ip2(\cache_data[5][20] ), .op(n9880) );
  nand4_1 U10086 ( .ip1(n9883), .ip2(n9882), .ip3(n9881), .ip4(n9880), .op(
        n9889) );
  nand2_1 U10087 ( .ip1(n12201), .ip2(\cache_data[4][20] ), .op(n9887) );
  nand2_1 U10088 ( .ip1(n12226), .ip2(\cache_data[7][20] ), .op(n9886) );
  nand2_1 U10089 ( .ip1(n12221), .ip2(\cache_data[15][20] ), .op(n9885) );
  nand2_1 U10090 ( .ip1(n12096), .ip2(\cache_data[11][20] ), .op(n9884) );
  nand4_1 U10091 ( .ip1(n9887), .ip2(n9886), .ip3(n9885), .ip4(n9884), .op(
        n9888) );
  or4_1 U10092 ( .ip1(n9891), .ip2(n9890), .ip3(n9889), .ip4(n9888), .op(
        n11193) );
  nand2_1 U10093 ( .ip1(n10828), .ip2(n11193), .op(n9956) );
  nand2_1 U10094 ( .ip1(n8894), .ip2(\cache_data[1][52] ), .op(n9895) );
  nand2_1 U10095 ( .ip1(n12219), .ip2(\cache_data[3][52] ), .op(n9894) );
  nand2_1 U10096 ( .ip1(n12241), .ip2(\cache_data[9][52] ), .op(n9893) );
  nand2_1 U10097 ( .ip1(n12233), .ip2(\cache_data[0][52] ), .op(n9892) );
  nand4_1 U10098 ( .ip1(n9895), .ip2(n9894), .ip3(n9893), .ip4(n9892), .op(
        n9911) );
  nand2_1 U10099 ( .ip1(n12202), .ip2(\cache_data[7][52] ), .op(n9899) );
  nand2_1 U10100 ( .ip1(n12191), .ip2(\cache_data[8][52] ), .op(n9898) );
  nand2_1 U10101 ( .ip1(n12179), .ip2(\cache_data[6][52] ), .op(n9897) );
  nand2_1 U10102 ( .ip1(n11927), .ip2(\cache_data[11][52] ), .op(n9896) );
  nand4_1 U10103 ( .ip1(n9899), .ip2(n9898), .ip3(n9897), .ip4(n9896), .op(
        n9910) );
  nand2_1 U10104 ( .ip1(n12235), .ip2(\cache_data[10][52] ), .op(n9903) );
  nand2_1 U10105 ( .ip1(n12220), .ip2(\cache_data[14][52] ), .op(n9902) );
  nand2_1 U10106 ( .ip1(n12228), .ip2(\cache_data[2][52] ), .op(n9901) );
  nand2_1 U10107 ( .ip1(n12243), .ip2(\cache_data[4][52] ), .op(n9900) );
  nand4_1 U10108 ( .ip1(n9903), .ip2(n9902), .ip3(n9901), .ip4(n9900), .op(
        n9909) );
  nand2_1 U10109 ( .ip1(n12165), .ip2(\cache_data[13][52] ), .op(n9907) );
  nand2_1 U10110 ( .ip1(n12221), .ip2(\cache_data[15][52] ), .op(n9906) );
  nand2_1 U10111 ( .ip1(n12240), .ip2(\cache_data[5][52] ), .op(n9905) );
  nand2_1 U10112 ( .ip1(n12227), .ip2(\cache_data[12][52] ), .op(n9904) );
  nand4_1 U10113 ( .ip1(n9907), .ip2(n9906), .ip3(n9905), .ip4(n9904), .op(
        n9908) );
  nor4_1 U10114 ( .ip1(n9911), .ip2(n9910), .ip3(n9909), .ip4(n9908), .op(
        n11194) );
  nor2_1 U10115 ( .ip1(n11194), .ip2(n10870), .op(n9933) );
  nand2_1 U10116 ( .ip1(n12165), .ip2(\cache_data[13][84] ), .op(n9915) );
  nand2_1 U10117 ( .ip1(n12221), .ip2(\cache_data[15][84] ), .op(n9914) );
  nand2_1 U10118 ( .ip1(n12233), .ip2(\cache_data[0][84] ), .op(n9913) );
  nand2_1 U10119 ( .ip1(n11927), .ip2(\cache_data[11][84] ), .op(n9912) );
  nand4_1 U10120 ( .ip1(n9915), .ip2(n9914), .ip3(n9913), .ip4(n9912), .op(
        n9931) );
  nand2_1 U10121 ( .ip1(n12228), .ip2(\cache_data[2][84] ), .op(n9919) );
  nand2_1 U10122 ( .ip1(n12179), .ip2(\cache_data[6][84] ), .op(n9918) );
  nand2_1 U10123 ( .ip1(n12191), .ip2(\cache_data[8][84] ), .op(n9917) );
  nand2_1 U10124 ( .ip1(n8894), .ip2(\cache_data[1][84] ), .op(n9916) );
  nand4_1 U10125 ( .ip1(n9919), .ip2(n9918), .ip3(n9917), .ip4(n9916), .op(
        n9930) );
  nand2_1 U10126 ( .ip1(n12219), .ip2(\cache_data[3][84] ), .op(n9923) );
  nand2_1 U10127 ( .ip1(n12235), .ip2(\cache_data[10][84] ), .op(n9922) );
  nand2_1 U10128 ( .ip1(n12220), .ip2(\cache_data[14][84] ), .op(n9921) );
  nand2_1 U10129 ( .ip1(n12240), .ip2(\cache_data[5][84] ), .op(n9920) );
  nand4_1 U10130 ( .ip1(n9923), .ip2(n9922), .ip3(n9921), .ip4(n9920), .op(
        n9929) );
  nand2_1 U10131 ( .ip1(n12243), .ip2(\cache_data[4][84] ), .op(n9927) );
  nand2_1 U10132 ( .ip1(n12227), .ip2(\cache_data[12][84] ), .op(n9926) );
  nand2_1 U10133 ( .ip1(n12241), .ip2(\cache_data[9][84] ), .op(n9925) );
  nand2_1 U10134 ( .ip1(n12202), .ip2(\cache_data[7][84] ), .op(n9924) );
  nand4_1 U10135 ( .ip1(n9927), .ip2(n9926), .ip3(n9925), .ip4(n9924), .op(
        n9928) );
  nor4_1 U10136 ( .ip1(n9931), .ip2(n9930), .ip3(n9929), .ip4(n9928), .op(
        n11195) );
  nor2_1 U10137 ( .ip1(n11195), .ip2(n10849), .op(n9932) );
  not_ab_or_c_or_d U10138 ( .ip1(data_wr_mem[20]), .ip2(n10873), .ip3(n9933), 
        .ip4(n9932), .op(n9955) );
  nand2_1 U10139 ( .ip1(n12179), .ip2(\cache_data[6][116] ), .op(n9937) );
  nand2_1 U10140 ( .ip1(n11943), .ip2(\cache_data[1][116] ), .op(n9936) );
  nand2_1 U10141 ( .ip1(n12096), .ip2(\cache_data[11][116] ), .op(n9935) );
  nand2_1 U10142 ( .ip1(n12207), .ip2(\cache_data[12][116] ), .op(n9934) );
  nand4_1 U10143 ( .ip1(n9937), .ip2(n9936), .ip3(n9935), .ip4(n9934), .op(
        n9953) );
  nand2_1 U10144 ( .ip1(n12240), .ip2(\cache_data[5][116] ), .op(n9941) );
  nand2_1 U10145 ( .ip1(n12235), .ip2(\cache_data[10][116] ), .op(n9940) );
  nand2_1 U10146 ( .ip1(n12233), .ip2(\cache_data[0][116] ), .op(n9939) );
  nand2_1 U10147 ( .ip1(n12201), .ip2(\cache_data[4][116] ), .op(n9938) );
  nand4_1 U10148 ( .ip1(n9941), .ip2(n9940), .ip3(n9939), .ip4(n9938), .op(
        n9952) );
  nand2_1 U10149 ( .ip1(n12142), .ip2(\cache_data[13][116] ), .op(n9945) );
  nand2_1 U10150 ( .ip1(n12126), .ip2(\cache_data[9][116] ), .op(n9944) );
  nand2_1 U10151 ( .ip1(n12121), .ip2(\cache_data[8][116] ), .op(n9943) );
  nand2_1 U10152 ( .ip1(n12219), .ip2(\cache_data[3][116] ), .op(n9942) );
  nand4_1 U10153 ( .ip1(n9945), .ip2(n9944), .ip3(n9943), .ip4(n9942), .op(
        n9951) );
  nand2_1 U10154 ( .ip1(n12226), .ip2(\cache_data[7][116] ), .op(n9949) );
  nand2_1 U10155 ( .ip1(n12221), .ip2(\cache_data[15][116] ), .op(n9948) );
  nand2_1 U10156 ( .ip1(n12220), .ip2(\cache_data[14][116] ), .op(n9947) );
  nand2_1 U10157 ( .ip1(n12228), .ip2(\cache_data[2][116] ), .op(n9946) );
  nand4_1 U10158 ( .ip1(n9949), .ip2(n9948), .ip3(n9947), .ip4(n9946), .op(
        n9950) );
  or4_1 U10159 ( .ip1(n9953), .ip2(n9952), .ip3(n9951), .ip4(n9950), .op(
        n11198) );
  nand2_1 U10160 ( .ip1(n10894), .ip2(n11198), .op(n9954) );
  nand3_1 U10161 ( .ip1(n9956), .ip2(n9955), .ip3(n9954), .op(n7428) );
  nand2_1 U10162 ( .ip1(data_wr_mem[21]), .ip2(n10873), .op(n10041) );
  nand2_1 U10163 ( .ip1(n12243), .ip2(\cache_data[4][117] ), .op(n9960) );
  nand2_1 U10164 ( .ip1(n12179), .ip2(\cache_data[6][117] ), .op(n9959) );
  nand2_1 U10165 ( .ip1(n8894), .ip2(\cache_data[1][117] ), .op(n9958) );
  nand2_1 U10166 ( .ip1(n12191), .ip2(\cache_data[8][117] ), .op(n9957) );
  nand4_1 U10167 ( .ip1(n9960), .ip2(n9959), .ip3(n9958), .ip4(n9957), .op(
        n9976) );
  nand2_1 U10168 ( .ip1(n11927), .ip2(\cache_data[11][117] ), .op(n9964) );
  nand2_1 U10169 ( .ip1(n9560), .ip2(\cache_data[12][117] ), .op(n9963) );
  nand2_1 U10170 ( .ip1(n12241), .ip2(\cache_data[9][117] ), .op(n9962) );
  nand2_1 U10171 ( .ip1(n12221), .ip2(\cache_data[15][117] ), .op(n9961) );
  nand4_1 U10172 ( .ip1(n9964), .ip2(n9963), .ip3(n9962), .ip4(n9961), .op(
        n9975) );
  nand2_1 U10173 ( .ip1(n12202), .ip2(\cache_data[7][117] ), .op(n9968) );
  nand2_1 U10174 ( .ip1(n12233), .ip2(\cache_data[0][117] ), .op(n9967) );
  nand2_1 U10175 ( .ip1(n12228), .ip2(\cache_data[2][117] ), .op(n9966) );
  nand2_1 U10176 ( .ip1(n12165), .ip2(\cache_data[13][117] ), .op(n9965) );
  nand4_1 U10177 ( .ip1(n9968), .ip2(n9967), .ip3(n9966), .ip4(n9965), .op(
        n9974) );
  nand2_1 U10178 ( .ip1(n12240), .ip2(\cache_data[5][117] ), .op(n9972) );
  nand2_1 U10179 ( .ip1(n12220), .ip2(\cache_data[14][117] ), .op(n9971) );
  nand2_1 U10180 ( .ip1(n12235), .ip2(\cache_data[10][117] ), .op(n9970) );
  nand2_1 U10181 ( .ip1(n12219), .ip2(\cache_data[3][117] ), .op(n9969) );
  nand4_1 U10182 ( .ip1(n9972), .ip2(n9971), .ip3(n9970), .ip4(n9969), .op(
        n9973) );
  or4_1 U10183 ( .ip1(n9976), .ip2(n9975), .ip3(n9974), .ip4(n9973), .op(
        n11202) );
  nand2_1 U10184 ( .ip1(n12240), .ip2(\cache_data[5][85] ), .op(n9980) );
  nand2_1 U10185 ( .ip1(n12221), .ip2(\cache_data[15][85] ), .op(n9979) );
  nand2_1 U10186 ( .ip1(n12191), .ip2(\cache_data[8][85] ), .op(n9978) );
  nand2_1 U10187 ( .ip1(n11927), .ip2(\cache_data[11][85] ), .op(n9977) );
  nand4_1 U10188 ( .ip1(n9980), .ip2(n9979), .ip3(n9978), .ip4(n9977), .op(
        n9996) );
  nand2_1 U10189 ( .ip1(n12202), .ip2(\cache_data[7][85] ), .op(n9984) );
  nand2_1 U10190 ( .ip1(n12220), .ip2(\cache_data[14][85] ), .op(n9983) );
  nand2_1 U10191 ( .ip1(n12179), .ip2(\cache_data[6][85] ), .op(n9982) );
  nand2_1 U10192 ( .ip1(n9560), .ip2(\cache_data[12][85] ), .op(n9981) );
  nand4_1 U10193 ( .ip1(n9984), .ip2(n9983), .ip3(n9982), .ip4(n9981), .op(
        n9995) );
  nand2_1 U10194 ( .ip1(n8894), .ip2(\cache_data[1][85] ), .op(n9988) );
  nand2_1 U10195 ( .ip1(n12228), .ip2(\cache_data[2][85] ), .op(n9987) );
  nand2_1 U10196 ( .ip1(n12233), .ip2(\cache_data[0][85] ), .op(n9986) );
  nand2_1 U10197 ( .ip1(n12241), .ip2(\cache_data[9][85] ), .op(n9985) );
  nand4_1 U10198 ( .ip1(n9988), .ip2(n9987), .ip3(n9986), .ip4(n9985), .op(
        n9994) );
  nand2_1 U10199 ( .ip1(n12235), .ip2(\cache_data[10][85] ), .op(n9992) );
  nand2_1 U10200 ( .ip1(n12219), .ip2(\cache_data[3][85] ), .op(n9991) );
  nand2_1 U10201 ( .ip1(n12165), .ip2(\cache_data[13][85] ), .op(n9990) );
  nand2_1 U10202 ( .ip1(n12243), .ip2(\cache_data[4][85] ), .op(n9989) );
  nand4_1 U10203 ( .ip1(n9992), .ip2(n9991), .ip3(n9990), .ip4(n9989), .op(
        n9993) );
  nor4_1 U10204 ( .ip1(n9996), .ip2(n9995), .ip3(n9994), .ip4(n9993), .op(
        n11204) );
  nor2_1 U10205 ( .ip1(n11204), .ip2(n10849), .op(n10018) );
  nand2_1 U10206 ( .ip1(n12165), .ip2(\cache_data[13][53] ), .op(n10000) );
  nand2_1 U10207 ( .ip1(n8905), .ip2(\cache_data[6][53] ), .op(n9999) );
  nand2_1 U10208 ( .ip1(n12233), .ip2(\cache_data[0][53] ), .op(n9998) );
  nand2_1 U10209 ( .ip1(n12243), .ip2(\cache_data[4][53] ), .op(n9997) );
  nand4_1 U10210 ( .ip1(n10000), .ip2(n9999), .ip3(n9998), .ip4(n9997), .op(
        n10016) );
  nand2_1 U10211 ( .ip1(n9560), .ip2(\cache_data[12][53] ), .op(n10004) );
  nand2_1 U10212 ( .ip1(n12220), .ip2(\cache_data[14][53] ), .op(n10003) );
  nand2_1 U10213 ( .ip1(n9669), .ip2(\cache_data[11][53] ), .op(n10002) );
  nand2_1 U10214 ( .ip1(n8894), .ip2(\cache_data[1][53] ), .op(n10001) );
  nand4_1 U10215 ( .ip1(n10004), .ip2(n10003), .ip3(n10002), .ip4(n10001), 
        .op(n10015) );
  nand2_1 U10216 ( .ip1(n12221), .ip2(\cache_data[15][53] ), .op(n10008) );
  nand2_1 U10217 ( .ip1(n12191), .ip2(\cache_data[8][53] ), .op(n10007) );
  nand2_1 U10218 ( .ip1(n12202), .ip2(\cache_data[7][53] ), .op(n10006) );
  nand2_1 U10219 ( .ip1(n12241), .ip2(\cache_data[9][53] ), .op(n10005) );
  nand4_1 U10220 ( .ip1(n10008), .ip2(n10007), .ip3(n10006), .ip4(n10005), 
        .op(n10014) );
  nand2_1 U10221 ( .ip1(n12219), .ip2(\cache_data[3][53] ), .op(n10012) );
  nand2_1 U10222 ( .ip1(n12196), .ip2(\cache_data[10][53] ), .op(n10011) );
  nand2_1 U10223 ( .ip1(n12240), .ip2(\cache_data[5][53] ), .op(n10010) );
  nand2_1 U10224 ( .ip1(n12228), .ip2(\cache_data[2][53] ), .op(n10009) );
  nand4_1 U10225 ( .ip1(n10012), .ip2(n10011), .ip3(n10010), .ip4(n10009), 
        .op(n10013) );
  nor4_1 U10226 ( .ip1(n10016), .ip2(n10015), .ip3(n10014), .ip4(n10013), .op(
        n11203) );
  nor2_1 U10227 ( .ip1(n11203), .ip2(n10870), .op(n10017) );
  not_ab_or_c_or_d U10228 ( .ip1(n10894), .ip2(n11202), .ip3(n10018), .ip4(
        n10017), .op(n10040) );
  nand2_1 U10229 ( .ip1(n12191), .ip2(\cache_data[8][21] ), .op(n10022) );
  nand2_1 U10230 ( .ip1(n12243), .ip2(\cache_data[4][21] ), .op(n10021) );
  nand2_1 U10231 ( .ip1(n12179), .ip2(\cache_data[6][21] ), .op(n10020) );
  nand2_1 U10232 ( .ip1(n12228), .ip2(\cache_data[2][21] ), .op(n10019) );
  nand4_1 U10233 ( .ip1(n10022), .ip2(n10021), .ip3(n10020), .ip4(n10019), 
        .op(n10038) );
  nand2_1 U10234 ( .ip1(n12202), .ip2(\cache_data[7][21] ), .op(n10026) );
  nand2_1 U10235 ( .ip1(n12240), .ip2(\cache_data[5][21] ), .op(n10025) );
  nand2_1 U10236 ( .ip1(n11927), .ip2(\cache_data[11][21] ), .op(n10024) );
  nand2_1 U10237 ( .ip1(n12165), .ip2(\cache_data[13][21] ), .op(n10023) );
  nand4_1 U10238 ( .ip1(n10026), .ip2(n10025), .ip3(n10024), .ip4(n10023), 
        .op(n10037) );
  nand2_1 U10239 ( .ip1(n12220), .ip2(\cache_data[14][21] ), .op(n10030) );
  nand2_1 U10240 ( .ip1(n12221), .ip2(\cache_data[15][21] ), .op(n10029) );
  nand2_1 U10241 ( .ip1(n8894), .ip2(\cache_data[1][21] ), .op(n10028) );
  nand2_1 U10242 ( .ip1(n12241), .ip2(\cache_data[9][21] ), .op(n10027) );
  nand4_1 U10243 ( .ip1(n10030), .ip2(n10029), .ip3(n10028), .ip4(n10027), 
        .op(n10036) );
  nand2_1 U10244 ( .ip1(n9560), .ip2(\cache_data[12][21] ), .op(n10034) );
  nand2_1 U10245 ( .ip1(n12219), .ip2(\cache_data[3][21] ), .op(n10033) );
  nand2_1 U10246 ( .ip1(n12233), .ip2(\cache_data[0][21] ), .op(n10032) );
  nand2_1 U10247 ( .ip1(n12235), .ip2(\cache_data[10][21] ), .op(n10031) );
  nand4_1 U10248 ( .ip1(n10034), .ip2(n10033), .ip3(n10032), .ip4(n10031), 
        .op(n10035) );
  or4_1 U10249 ( .ip1(n10038), .ip2(n10037), .ip3(n10036), .ip4(n10035), .op(
        n11207) );
  nand2_1 U10250 ( .ip1(n10828), .ip2(n11207), .op(n10039) );
  nand3_1 U10251 ( .ip1(n10041), .ip2(n10040), .ip3(n10039), .op(n7427) );
  nand2_1 U10252 ( .ip1(n12228), .ip2(\cache_data[2][22] ), .op(n10045) );
  nand2_1 U10253 ( .ip1(n12240), .ip2(\cache_data[5][22] ), .op(n10044) );
  nand2_1 U10254 ( .ip1(n12207), .ip2(\cache_data[12][22] ), .op(n10043) );
  nand2_1 U10255 ( .ip1(n12121), .ip2(\cache_data[8][22] ), .op(n10042) );
  nand4_1 U10256 ( .ip1(n10045), .ip2(n10044), .ip3(n10043), .ip4(n10042), 
        .op(n10061) );
  nand2_1 U10257 ( .ip1(n12126), .ip2(\cache_data[9][22] ), .op(n10049) );
  nand2_1 U10258 ( .ip1(n12226), .ip2(\cache_data[7][22] ), .op(n10048) );
  nand2_1 U10259 ( .ip1(n12196), .ip2(\cache_data[10][22] ), .op(n10047) );
  nand2_1 U10260 ( .ip1(n12221), .ip2(\cache_data[15][22] ), .op(n10046) );
  nand4_1 U10261 ( .ip1(n10049), .ip2(n10048), .ip3(n10047), .ip4(n10046), 
        .op(n10060) );
  nand2_1 U10262 ( .ip1(n12219), .ip2(\cache_data[3][22] ), .op(n10053) );
  nand2_1 U10263 ( .ip1(n12201), .ip2(\cache_data[4][22] ), .op(n10052) );
  nand2_1 U10264 ( .ip1(n12233), .ip2(\cache_data[0][22] ), .op(n10051) );
  nand2_1 U10265 ( .ip1(n10305), .ip2(\cache_data[6][22] ), .op(n10050) );
  nand4_1 U10266 ( .ip1(n10053), .ip2(n10052), .ip3(n10051), .ip4(n10050), 
        .op(n10059) );
  nand2_1 U10267 ( .ip1(n12220), .ip2(\cache_data[14][22] ), .op(n10057) );
  nand2_1 U10268 ( .ip1(n11979), .ip2(\cache_data[1][22] ), .op(n10056) );
  nand2_1 U10269 ( .ip1(n9669), .ip2(\cache_data[11][22] ), .op(n10055) );
  nand2_1 U10270 ( .ip1(n12142), .ip2(\cache_data[13][22] ), .op(n10054) );
  nand4_1 U10271 ( .ip1(n10057), .ip2(n10056), .ip3(n10055), .ip4(n10054), 
        .op(n10058) );
  or4_1 U10272 ( .ip1(n10061), .ip2(n10060), .ip3(n10059), .ip4(n10058), .op(
        n11216) );
  nand2_1 U10273 ( .ip1(n10828), .ip2(n11216), .op(n10126) );
  nand2_1 U10274 ( .ip1(n9669), .ip2(\cache_data[11][54] ), .op(n10065) );
  nand2_1 U10275 ( .ip1(n12196), .ip2(\cache_data[10][54] ), .op(n10064) );
  nand2_1 U10276 ( .ip1(n12221), .ip2(\cache_data[15][54] ), .op(n10063) );
  nand2_1 U10277 ( .ip1(n12165), .ip2(\cache_data[13][54] ), .op(n10062) );
  nand4_1 U10278 ( .ip1(n10065), .ip2(n10064), .ip3(n10063), .ip4(n10062), 
        .op(n10081) );
  nand2_1 U10279 ( .ip1(n12219), .ip2(\cache_data[3][54] ), .op(n10069) );
  nand2_1 U10280 ( .ip1(n12241), .ip2(\cache_data[9][54] ), .op(n10068) );
  nand2_1 U10281 ( .ip1(n12191), .ip2(\cache_data[8][54] ), .op(n10067) );
  nand2_1 U10282 ( .ip1(n12233), .ip2(\cache_data[0][54] ), .op(n10066) );
  nand4_1 U10283 ( .ip1(n10069), .ip2(n10068), .ip3(n10067), .ip4(n10066), 
        .op(n10080) );
  nand2_1 U10284 ( .ip1(n12243), .ip2(\cache_data[4][54] ), .op(n10073) );
  nand2_1 U10285 ( .ip1(n8894), .ip2(\cache_data[1][54] ), .op(n10072) );
  nand2_1 U10286 ( .ip1(n12202), .ip2(\cache_data[7][54] ), .op(n10071) );
  nand2_1 U10287 ( .ip1(n12228), .ip2(\cache_data[2][54] ), .op(n10070) );
  nand4_1 U10288 ( .ip1(n10073), .ip2(n10072), .ip3(n10071), .ip4(n10070), 
        .op(n10079) );
  nand2_1 U10289 ( .ip1(n8905), .ip2(\cache_data[6][54] ), .op(n10077) );
  nand2_1 U10290 ( .ip1(n9560), .ip2(\cache_data[12][54] ), .op(n10076) );
  nand2_1 U10291 ( .ip1(n12240), .ip2(\cache_data[5][54] ), .op(n10075) );
  nand2_1 U10292 ( .ip1(n12220), .ip2(\cache_data[14][54] ), .op(n10074) );
  nand4_1 U10293 ( .ip1(n10077), .ip2(n10076), .ip3(n10075), .ip4(n10074), 
        .op(n10078) );
  nor4_1 U10294 ( .ip1(n10081), .ip2(n10080), .ip3(n10079), .ip4(n10078), .op(
        n11213) );
  nor2_1 U10295 ( .ip1(n11213), .ip2(n10870), .op(n10103) );
  nand2_1 U10296 ( .ip1(n12219), .ip2(\cache_data[3][86] ), .op(n10085) );
  nand2_1 U10297 ( .ip1(n12165), .ip2(\cache_data[13][86] ), .op(n10084) );
  nand2_1 U10298 ( .ip1(n12191), .ip2(\cache_data[8][86] ), .op(n10083) );
  nand2_1 U10299 ( .ip1(n12241), .ip2(\cache_data[9][86] ), .op(n10082) );
  nand4_1 U10300 ( .ip1(n10085), .ip2(n10084), .ip3(n10083), .ip4(n10082), 
        .op(n10101) );
  nand2_1 U10301 ( .ip1(n12233), .ip2(\cache_data[0][86] ), .op(n10089) );
  nand2_1 U10302 ( .ip1(n12202), .ip2(\cache_data[7][86] ), .op(n10088) );
  nand2_1 U10303 ( .ip1(n12243), .ip2(\cache_data[4][86] ), .op(n10087) );
  nand2_1 U10304 ( .ip1(n11927), .ip2(\cache_data[11][86] ), .op(n10086) );
  nand4_1 U10305 ( .ip1(n10089), .ip2(n10088), .ip3(n10087), .ip4(n10086), 
        .op(n10100) );
  nand2_1 U10306 ( .ip1(n8894), .ip2(\cache_data[1][86] ), .op(n10093) );
  nand2_1 U10307 ( .ip1(n12227), .ip2(\cache_data[12][86] ), .op(n10092) );
  nand2_1 U10308 ( .ip1(n12240), .ip2(\cache_data[5][86] ), .op(n10091) );
  nand2_1 U10309 ( .ip1(n12179), .ip2(\cache_data[6][86] ), .op(n10090) );
  nand4_1 U10310 ( .ip1(n10093), .ip2(n10092), .ip3(n10091), .ip4(n10090), 
        .op(n10099) );
  nand2_1 U10311 ( .ip1(n12221), .ip2(\cache_data[15][86] ), .op(n10097) );
  nand2_1 U10312 ( .ip1(n12220), .ip2(\cache_data[14][86] ), .op(n10096) );
  nand2_1 U10313 ( .ip1(n12228), .ip2(\cache_data[2][86] ), .op(n10095) );
  nand2_1 U10314 ( .ip1(n12235), .ip2(\cache_data[10][86] ), .op(n10094) );
  nand4_1 U10315 ( .ip1(n10097), .ip2(n10096), .ip3(n10095), .ip4(n10094), 
        .op(n10098) );
  nor4_1 U10316 ( .ip1(n10101), .ip2(n10100), .ip3(n10099), .ip4(n10098), .op(
        n11212) );
  nor2_1 U10317 ( .ip1(n11212), .ip2(n10849), .op(n10102) );
  not_ab_or_c_or_d U10318 ( .ip1(data_wr_mem[22]), .ip2(n10873), .ip3(n10103), 
        .ip4(n10102), .op(n10125) );
  nand2_1 U10319 ( .ip1(n12226), .ip2(\cache_data[7][118] ), .op(n10107) );
  nand2_1 U10320 ( .ip1(n12121), .ip2(\cache_data[8][118] ), .op(n10106) );
  nand2_1 U10321 ( .ip1(n10305), .ip2(\cache_data[6][118] ), .op(n10105) );
  nand2_1 U10322 ( .ip1(n12142), .ip2(\cache_data[13][118] ), .op(n10104) );
  nand4_1 U10323 ( .ip1(n10107), .ip2(n10106), .ip3(n10105), .ip4(n10104), 
        .op(n10123) );
  nand2_1 U10324 ( .ip1(n12228), .ip2(\cache_data[2][118] ), .op(n10111) );
  nand2_1 U10325 ( .ip1(n12240), .ip2(\cache_data[5][118] ), .op(n10110) );
  nand2_1 U10326 ( .ip1(n12207), .ip2(\cache_data[12][118] ), .op(n10109) );
  nand2_1 U10327 ( .ip1(n9669), .ip2(\cache_data[11][118] ), .op(n10108) );
  nand4_1 U10328 ( .ip1(n10111), .ip2(n10110), .ip3(n10109), .ip4(n10108), 
        .op(n10122) );
  nand2_1 U10329 ( .ip1(n12233), .ip2(\cache_data[0][118] ), .op(n10115) );
  nand2_1 U10330 ( .ip1(n11943), .ip2(\cache_data[1][118] ), .op(n10114) );
  nand2_1 U10331 ( .ip1(n12126), .ip2(\cache_data[9][118] ), .op(n10113) );
  nand2_1 U10332 ( .ip1(n12221), .ip2(\cache_data[15][118] ), .op(n10112) );
  nand4_1 U10333 ( .ip1(n10115), .ip2(n10114), .ip3(n10113), .ip4(n10112), 
        .op(n10121) );
  nand2_1 U10334 ( .ip1(n12219), .ip2(\cache_data[3][118] ), .op(n10119) );
  nand2_1 U10335 ( .ip1(n12196), .ip2(\cache_data[10][118] ), .op(n10118) );
  nand2_1 U10336 ( .ip1(n12201), .ip2(\cache_data[4][118] ), .op(n10117) );
  nand2_1 U10337 ( .ip1(n12220), .ip2(\cache_data[14][118] ), .op(n10116) );
  nand4_1 U10338 ( .ip1(n10119), .ip2(n10118), .ip3(n10117), .ip4(n10116), 
        .op(n10120) );
  or4_1 U10339 ( .ip1(n10123), .ip2(n10122), .ip3(n10121), .ip4(n10120), .op(
        n11211) );
  nand2_1 U10340 ( .ip1(n10894), .ip2(n11211), .op(n10124) );
  nand3_1 U10341 ( .ip1(n10126), .ip2(n10125), .ip3(n10124), .op(n7426) );
  nand2_1 U10342 ( .ip1(n12228), .ip2(\cache_data[2][23] ), .op(n10130) );
  nand2_1 U10343 ( .ip1(n12221), .ip2(\cache_data[15][23] ), .op(n10129) );
  nand2_1 U10344 ( .ip1(n9560), .ip2(\cache_data[12][23] ), .op(n10128) );
  nand2_1 U10345 ( .ip1(n10305), .ip2(\cache_data[6][23] ), .op(n10127) );
  nand4_1 U10346 ( .ip1(n10130), .ip2(n10129), .ip3(n10128), .ip4(n10127), 
        .op(n10146) );
  nand2_1 U10347 ( .ip1(n12220), .ip2(\cache_data[14][23] ), .op(n10134) );
  nand2_1 U10348 ( .ip1(n12191), .ip2(\cache_data[8][23] ), .op(n10133) );
  nand2_1 U10349 ( .ip1(n8894), .ip2(\cache_data[1][23] ), .op(n10132) );
  nand2_1 U10350 ( .ip1(n9669), .ip2(\cache_data[11][23] ), .op(n10131) );
  nand4_1 U10351 ( .ip1(n10134), .ip2(n10133), .ip3(n10132), .ip4(n10131), 
        .op(n10145) );
  nand2_1 U10352 ( .ip1(n12240), .ip2(\cache_data[5][23] ), .op(n10138) );
  nand2_1 U10353 ( .ip1(n12165), .ip2(\cache_data[13][23] ), .op(n10137) );
  nand2_1 U10354 ( .ip1(n12233), .ip2(\cache_data[0][23] ), .op(n10136) );
  nand2_1 U10355 ( .ip1(n12241), .ip2(\cache_data[9][23] ), .op(n10135) );
  nand4_1 U10356 ( .ip1(n10138), .ip2(n10137), .ip3(n10136), .ip4(n10135), 
        .op(n10144) );
  nand2_1 U10357 ( .ip1(n12196), .ip2(\cache_data[10][23] ), .op(n10142) );
  nand2_1 U10358 ( .ip1(n12202), .ip2(\cache_data[7][23] ), .op(n10141) );
  nand2_1 U10359 ( .ip1(n12219), .ip2(\cache_data[3][23] ), .op(n10140) );
  nand2_1 U10360 ( .ip1(n12243), .ip2(\cache_data[4][23] ), .op(n10139) );
  nand4_1 U10361 ( .ip1(n10142), .ip2(n10141), .ip3(n10140), .ip4(n10139), 
        .op(n10143) );
  or4_1 U10362 ( .ip1(n10146), .ip2(n10145), .ip3(n10144), .ip4(n10143), .op(
        n11225) );
  nand2_1 U10363 ( .ip1(n10828), .ip2(n11225), .op(n10211) );
  nand2_1 U10364 ( .ip1(n11927), .ip2(\cache_data[11][55] ), .op(n10150) );
  nand2_1 U10365 ( .ip1(n12202), .ip2(\cache_data[7][55] ), .op(n10149) );
  nand2_1 U10366 ( .ip1(n12219), .ip2(\cache_data[3][55] ), .op(n10148) );
  nand2_1 U10367 ( .ip1(n12191), .ip2(\cache_data[8][55] ), .op(n10147) );
  nand4_1 U10368 ( .ip1(n10150), .ip2(n10149), .ip3(n10148), .ip4(n10147), 
        .op(n10166) );
  nand2_1 U10369 ( .ip1(n12221), .ip2(\cache_data[15][55] ), .op(n10154) );
  nand2_1 U10370 ( .ip1(n12233), .ip2(\cache_data[0][55] ), .op(n10153) );
  nand2_1 U10371 ( .ip1(n12227), .ip2(\cache_data[12][55] ), .op(n10152) );
  nand2_1 U10372 ( .ip1(n12240), .ip2(\cache_data[5][55] ), .op(n10151) );
  nand4_1 U10373 ( .ip1(n10154), .ip2(n10153), .ip3(n10152), .ip4(n10151), 
        .op(n10165) );
  nand2_1 U10374 ( .ip1(n12165), .ip2(\cache_data[13][55] ), .op(n10158) );
  nand2_1 U10375 ( .ip1(n12228), .ip2(\cache_data[2][55] ), .op(n10157) );
  nand2_1 U10376 ( .ip1(n12220), .ip2(\cache_data[14][55] ), .op(n10156) );
  nand2_1 U10377 ( .ip1(n12243), .ip2(\cache_data[4][55] ), .op(n10155) );
  nand4_1 U10378 ( .ip1(n10158), .ip2(n10157), .ip3(n10156), .ip4(n10155), 
        .op(n10164) );
  nand2_1 U10379 ( .ip1(n12179), .ip2(\cache_data[6][55] ), .op(n10162) );
  nand2_1 U10380 ( .ip1(n12241), .ip2(\cache_data[9][55] ), .op(n10161) );
  nand2_1 U10381 ( .ip1(n8894), .ip2(\cache_data[1][55] ), .op(n10160) );
  nand2_1 U10382 ( .ip1(n12235), .ip2(\cache_data[10][55] ), .op(n10159) );
  nand4_1 U10383 ( .ip1(n10162), .ip2(n10161), .ip3(n10160), .ip4(n10159), 
        .op(n10163) );
  nor4_1 U10384 ( .ip1(n10166), .ip2(n10165), .ip3(n10164), .ip4(n10163), .op(
        n11222) );
  nor2_1 U10385 ( .ip1(n11222), .ip2(n10870), .op(n10188) );
  nand2_1 U10386 ( .ip1(n12165), .ip2(\cache_data[13][87] ), .op(n10170) );
  nand2_1 U10387 ( .ip1(n12191), .ip2(\cache_data[8][87] ), .op(n10169) );
  nand2_1 U10388 ( .ip1(n12219), .ip2(\cache_data[3][87] ), .op(n10168) );
  nand2_1 U10389 ( .ip1(n8894), .ip2(\cache_data[1][87] ), .op(n10167) );
  nand4_1 U10390 ( .ip1(n10170), .ip2(n10169), .ip3(n10168), .ip4(n10167), 
        .op(n10186) );
  nand2_1 U10391 ( .ip1(n12241), .ip2(\cache_data[9][87] ), .op(n10174) );
  nand2_1 U10392 ( .ip1(n12220), .ip2(\cache_data[14][87] ), .op(n10173) );
  nand2_1 U10393 ( .ip1(n12196), .ip2(\cache_data[10][87] ), .op(n10172) );
  nand2_1 U10394 ( .ip1(n12221), .ip2(\cache_data[15][87] ), .op(n10171) );
  nand4_1 U10395 ( .ip1(n10174), .ip2(n10173), .ip3(n10172), .ip4(n10171), 
        .op(n10185) );
  nand2_1 U10396 ( .ip1(n9669), .ip2(\cache_data[11][87] ), .op(n10178) );
  nand2_1 U10397 ( .ip1(n12202), .ip2(\cache_data[7][87] ), .op(n10177) );
  nand2_1 U10398 ( .ip1(n12240), .ip2(\cache_data[5][87] ), .op(n10176) );
  nand2_1 U10399 ( .ip1(n12233), .ip2(\cache_data[0][87] ), .op(n10175) );
  nand4_1 U10400 ( .ip1(n10178), .ip2(n10177), .ip3(n10176), .ip4(n10175), 
        .op(n10184) );
  nand2_1 U10401 ( .ip1(n12228), .ip2(\cache_data[2][87] ), .op(n10182) );
  nand2_1 U10402 ( .ip1(n12227), .ip2(\cache_data[12][87] ), .op(n10181) );
  nand2_1 U10403 ( .ip1(n8905), .ip2(\cache_data[6][87] ), .op(n10180) );
  nand2_1 U10404 ( .ip1(n12243), .ip2(\cache_data[4][87] ), .op(n10179) );
  nand4_1 U10405 ( .ip1(n10182), .ip2(n10181), .ip3(n10180), .ip4(n10179), 
        .op(n10183) );
  nor4_1 U10406 ( .ip1(n10186), .ip2(n10185), .ip3(n10184), .ip4(n10183), .op(
        n11221) );
  nor2_1 U10407 ( .ip1(n11221), .ip2(n10849), .op(n10187) );
  not_ab_or_c_or_d U10408 ( .ip1(data_wr_mem[23]), .ip2(n10873), .ip3(n10188), 
        .ip4(n10187), .op(n10210) );
  nand2_1 U10409 ( .ip1(n12226), .ip2(\cache_data[7][119] ), .op(n10192) );
  nand2_1 U10410 ( .ip1(n10305), .ip2(\cache_data[6][119] ), .op(n10191) );
  nand2_1 U10411 ( .ip1(n9560), .ip2(\cache_data[12][119] ), .op(n10190) );
  nand2_1 U10412 ( .ip1(n12121), .ip2(\cache_data[8][119] ), .op(n10189) );
  nand4_1 U10413 ( .ip1(n10192), .ip2(n10191), .ip3(n10190), .ip4(n10189), 
        .op(n10208) );
  nand2_1 U10414 ( .ip1(n12221), .ip2(\cache_data[15][119] ), .op(n10196) );
  nand2_1 U10415 ( .ip1(n9669), .ip2(\cache_data[11][119] ), .op(n10195) );
  nand2_1 U10416 ( .ip1(n12126), .ip2(\cache_data[9][119] ), .op(n10194) );
  nand2_1 U10417 ( .ip1(n12228), .ip2(\cache_data[2][119] ), .op(n10193) );
  nand4_1 U10418 ( .ip1(n10196), .ip2(n10195), .ip3(n10194), .ip4(n10193), 
        .op(n10207) );
  nand2_1 U10419 ( .ip1(n12196), .ip2(\cache_data[10][119] ), .op(n10200) );
  nand2_1 U10420 ( .ip1(n12201), .ip2(\cache_data[4][119] ), .op(n10199) );
  nand2_1 U10421 ( .ip1(n12220), .ip2(\cache_data[14][119] ), .op(n10198) );
  nand2_1 U10422 ( .ip1(n12219), .ip2(\cache_data[3][119] ), .op(n10197) );
  nand4_1 U10423 ( .ip1(n10200), .ip2(n10199), .ip3(n10198), .ip4(n10197), 
        .op(n10206) );
  nand2_1 U10424 ( .ip1(n12233), .ip2(\cache_data[0][119] ), .op(n10204) );
  nand2_1 U10425 ( .ip1(n12142), .ip2(\cache_data[13][119] ), .op(n10203) );
  nand2_1 U10426 ( .ip1(n11979), .ip2(\cache_data[1][119] ), .op(n10202) );
  nand2_1 U10427 ( .ip1(n12240), .ip2(\cache_data[5][119] ), .op(n10201) );
  nand4_1 U10428 ( .ip1(n10204), .ip2(n10203), .ip3(n10202), .ip4(n10201), 
        .op(n10205) );
  or4_1 U10429 ( .ip1(n10208), .ip2(n10207), .ip3(n10206), .ip4(n10205), .op(
        n11220) );
  nand2_1 U10430 ( .ip1(n10894), .ip2(n11220), .op(n10209) );
  nand3_1 U10431 ( .ip1(n10211), .ip2(n10210), .ip3(n10209), .op(n7425) );
  nand2_1 U10432 ( .ip1(n12227), .ip2(\cache_data[12][24] ), .op(n10215) );
  inv_1 U10433 ( .ip(n8928), .op(n11973) );
  nand2_1 U10434 ( .ip1(n11973), .ip2(\cache_data[2][24] ), .op(n10214) );
  nand2_1 U10435 ( .ip1(n12152), .ip2(\cache_data[9][24] ), .op(n10213) );
  nand2_1 U10436 ( .ip1(n12165), .ip2(\cache_data[13][24] ), .op(n10212) );
  nand4_1 U10437 ( .ip1(n10215), .ip2(n10214), .ip3(n10213), .ip4(n10212), 
        .op(n10231) );
  inv_1 U10438 ( .ip(n8923), .op(n11964) );
  nand2_1 U10439 ( .ip1(n11964), .ip2(\cache_data[0][24] ), .op(n10219) );
  inv_1 U10440 ( .ip(n8146), .op(n11966) );
  nand2_1 U10441 ( .ip1(n11966), .ip2(\cache_data[10][24] ), .op(n10218) );
  inv_1 U10442 ( .ip(n10964), .op(n11493) );
  inv_1 U10443 ( .ip(n11493), .op(n11963) );
  nand2_1 U10444 ( .ip1(n11963), .ip2(\cache_data[5][24] ), .op(n10217) );
  inv_1 U10445 ( .ip(n10975), .op(n11612) );
  inv_1 U10446 ( .ip(n11612), .op(n11965) );
  nand2_1 U10447 ( .ip1(n11965), .ip2(\cache_data[15][24] ), .op(n10216) );
  nand4_1 U10448 ( .ip1(n10219), .ip2(n10218), .ip3(n10217), .ip4(n10216), 
        .op(n10230) );
  nand2_1 U10449 ( .ip1(n12164), .ip2(\cache_data[4][24] ), .op(n10223) );
  inv_1 U10450 ( .ip(n10305), .op(n11502) );
  inv_1 U10451 ( .ip(n11502), .op(n11972) );
  nand2_1 U10452 ( .ip1(n11972), .ip2(\cache_data[6][24] ), .op(n10222) );
  nand2_1 U10453 ( .ip1(n12191), .ip2(\cache_data[8][24] ), .op(n10221) );
  inv_1 U10454 ( .ip(n12120), .op(n11459) );
  inv_1 U10455 ( .ip(n11459), .op(n11943) );
  nand2_1 U10456 ( .ip1(n11943), .ip2(\cache_data[1][24] ), .op(n10220) );
  nand4_1 U10457 ( .ip1(n10223), .ip2(n10222), .ip3(n10221), .ip4(n10220), 
        .op(n10229) );
  nand2_1 U10458 ( .ip1(n12143), .ip2(\cache_data[7][24] ), .op(n10227) );
  nand2_1 U10459 ( .ip1(n11688), .ip2(\cache_data[14][24] ), .op(n10226) );
  inv_1 U10460 ( .ip(n12219), .op(n11476) );
  inv_1 U10461 ( .ip(n11476), .op(n11978) );
  nand2_1 U10462 ( .ip1(n11978), .ip2(\cache_data[3][24] ), .op(n10225) );
  nand2_1 U10463 ( .ip1(n11927), .ip2(\cache_data[11][24] ), .op(n10224) );
  nand4_1 U10464 ( .ip1(n10227), .ip2(n10226), .ip3(n10225), .ip4(n10224), 
        .op(n10228) );
  or4_1 U10465 ( .ip1(n10231), .ip2(n10230), .ip3(n10229), .ip4(n10228), .op(
        n11229) );
  nand2_1 U10466 ( .ip1(n10828), .ip2(n11229), .op(n10296) );
  nand2_1 U10467 ( .ip1(n11964), .ip2(\cache_data[0][56] ), .op(n10235) );
  nand2_1 U10468 ( .ip1(n11943), .ip2(\cache_data[1][56] ), .op(n10234) );
  nand2_1 U10469 ( .ip1(n12143), .ip2(\cache_data[7][56] ), .op(n10233) );
  nand2_1 U10470 ( .ip1(n12191), .ip2(\cache_data[8][56] ), .op(n10232) );
  nand4_1 U10471 ( .ip1(n10235), .ip2(n10234), .ip3(n10233), .ip4(n10232), 
        .op(n10251) );
  nand2_1 U10472 ( .ip1(n11963), .ip2(\cache_data[5][56] ), .op(n10239) );
  nand2_1 U10473 ( .ip1(n12227), .ip2(\cache_data[12][56] ), .op(n10238) );
  nand2_1 U10474 ( .ip1(n12164), .ip2(\cache_data[4][56] ), .op(n10237) );
  nand2_1 U10475 ( .ip1(n11972), .ip2(\cache_data[6][56] ), .op(n10236) );
  nand4_1 U10476 ( .ip1(n10239), .ip2(n10238), .ip3(n10237), .ip4(n10236), 
        .op(n10250) );
  nand2_1 U10477 ( .ip1(n11978), .ip2(\cache_data[3][56] ), .op(n10243) );
  nand2_1 U10478 ( .ip1(n11927), .ip2(\cache_data[11][56] ), .op(n10242) );
  nand2_1 U10479 ( .ip1(n12152), .ip2(\cache_data[9][56] ), .op(n10241) );
  nand2_1 U10480 ( .ip1(n12165), .ip2(\cache_data[13][56] ), .op(n10240) );
  nand4_1 U10481 ( .ip1(n10243), .ip2(n10242), .ip3(n10241), .ip4(n10240), 
        .op(n10249) );
  nand2_1 U10482 ( .ip1(n11965), .ip2(\cache_data[15][56] ), .op(n10247) );
  nand2_1 U10483 ( .ip1(n11966), .ip2(\cache_data[10][56] ), .op(n10246) );
  nand2_1 U10484 ( .ip1(n11688), .ip2(\cache_data[14][56] ), .op(n10245) );
  nand2_1 U10485 ( .ip1(n11973), .ip2(\cache_data[2][56] ), .op(n10244) );
  nand4_1 U10486 ( .ip1(n10247), .ip2(n10246), .ip3(n10245), .ip4(n10244), 
        .op(n10248) );
  nor4_1 U10487 ( .ip1(n10251), .ip2(n10250), .ip3(n10249), .ip4(n10248), .op(
        n11231) );
  nor2_1 U10488 ( .ip1(n11231), .ip2(n10870), .op(n10273) );
  nand2_1 U10489 ( .ip1(n11963), .ip2(\cache_data[5][88] ), .op(n10255) );
  nand2_1 U10490 ( .ip1(n11688), .ip2(\cache_data[14][88] ), .op(n10254) );
  nand2_1 U10491 ( .ip1(n11943), .ip2(\cache_data[1][88] ), .op(n10253) );
  nand2_1 U10492 ( .ip1(n12191), .ip2(\cache_data[8][88] ), .op(n10252) );
  nand4_1 U10493 ( .ip1(n10255), .ip2(n10254), .ip3(n10253), .ip4(n10252), 
        .op(n10271) );
  nand2_1 U10494 ( .ip1(n12164), .ip2(\cache_data[4][88] ), .op(n10259) );
  nand2_1 U10495 ( .ip1(n12152), .ip2(\cache_data[9][88] ), .op(n10258) );
  nand2_1 U10496 ( .ip1(n11966), .ip2(\cache_data[10][88] ), .op(n10257) );
  nand2_1 U10497 ( .ip1(n11965), .ip2(\cache_data[15][88] ), .op(n10256) );
  nand4_1 U10498 ( .ip1(n10259), .ip2(n10258), .ip3(n10257), .ip4(n10256), 
        .op(n10270) );
  nand2_1 U10499 ( .ip1(n12165), .ip2(\cache_data[13][88] ), .op(n10263) );
  nand2_1 U10500 ( .ip1(n11927), .ip2(\cache_data[11][88] ), .op(n10262) );
  nand2_1 U10501 ( .ip1(n11964), .ip2(\cache_data[0][88] ), .op(n10261) );
  nand2_1 U10502 ( .ip1(n11973), .ip2(\cache_data[2][88] ), .op(n10260) );
  nand4_1 U10503 ( .ip1(n10263), .ip2(n10262), .ip3(n10261), .ip4(n10260), 
        .op(n10269) );
  nand2_1 U10504 ( .ip1(n12143), .ip2(\cache_data[7][88] ), .op(n10267) );
  nand2_1 U10505 ( .ip1(n12227), .ip2(\cache_data[12][88] ), .op(n10266) );
  nand2_1 U10506 ( .ip1(n11978), .ip2(\cache_data[3][88] ), .op(n10265) );
  nand2_1 U10507 ( .ip1(n11972), .ip2(\cache_data[6][88] ), .op(n10264) );
  nand4_1 U10508 ( .ip1(n10267), .ip2(n10266), .ip3(n10265), .ip4(n10264), 
        .op(n10268) );
  nor4_1 U10509 ( .ip1(n10271), .ip2(n10270), .ip3(n10269), .ip4(n10268), .op(
        n11230) );
  nor2_1 U10510 ( .ip1(n11230), .ip2(n10849), .op(n10272) );
  not_ab_or_c_or_d U10511 ( .ip1(data_wr_mem[24]), .ip2(n10873), .ip3(n10273), 
        .ip4(n10272), .op(n10295) );
  nand2_1 U10512 ( .ip1(n11943), .ip2(\cache_data[1][120] ), .op(n10277) );
  nand2_1 U10513 ( .ip1(n11965), .ip2(\cache_data[15][120] ), .op(n10276) );
  nand2_1 U10514 ( .ip1(n11978), .ip2(\cache_data[3][120] ), .op(n10275) );
  nand2_1 U10515 ( .ip1(n12191), .ip2(\cache_data[8][120] ), .op(n10274) );
  nand4_1 U10516 ( .ip1(n10277), .ip2(n10276), .ip3(n10275), .ip4(n10274), 
        .op(n10293) );
  nand2_1 U10517 ( .ip1(n12152), .ip2(\cache_data[9][120] ), .op(n10281) );
  nand2_1 U10518 ( .ip1(n11964), .ip2(\cache_data[0][120] ), .op(n10280) );
  nand2_1 U10519 ( .ip1(n11688), .ip2(\cache_data[14][120] ), .op(n10279) );
  nand2_1 U10520 ( .ip1(n12164), .ip2(\cache_data[4][120] ), .op(n10278) );
  nand4_1 U10521 ( .ip1(n10281), .ip2(n10280), .ip3(n10279), .ip4(n10278), 
        .op(n10292) );
  nand2_1 U10522 ( .ip1(n11972), .ip2(\cache_data[6][120] ), .op(n10285) );
  nand2_1 U10523 ( .ip1(n11966), .ip2(\cache_data[10][120] ), .op(n10284) );
  nand2_1 U10524 ( .ip1(n12165), .ip2(\cache_data[13][120] ), .op(n10283) );
  nand2_1 U10525 ( .ip1(n12227), .ip2(\cache_data[12][120] ), .op(n10282) );
  nand4_1 U10526 ( .ip1(n10285), .ip2(n10284), .ip3(n10283), .ip4(n10282), 
        .op(n10291) );
  nand2_1 U10527 ( .ip1(n12143), .ip2(\cache_data[7][120] ), .op(n10289) );
  nand2_1 U10528 ( .ip1(n11973), .ip2(\cache_data[2][120] ), .op(n10288) );
  nand2_1 U10529 ( .ip1(n11963), .ip2(\cache_data[5][120] ), .op(n10287) );
  nand2_1 U10530 ( .ip1(n11927), .ip2(\cache_data[11][120] ), .op(n10286) );
  nand4_1 U10531 ( .ip1(n10289), .ip2(n10288), .ip3(n10287), .ip4(n10286), 
        .op(n10290) );
  or4_1 U10532 ( .ip1(n10293), .ip2(n10292), .ip3(n10291), .ip4(n10290), .op(
        n11234) );
  nand2_1 U10533 ( .ip1(n10894), .ip2(n11234), .op(n10294) );
  nand3_1 U10534 ( .ip1(n10296), .ip2(n10295), .ip3(n10294), .op(n7424) );
  nand2_1 U10535 ( .ip1(n12227), .ip2(\cache_data[12][25] ), .op(n10300) );
  nand2_1 U10536 ( .ip1(n12165), .ip2(\cache_data[13][25] ), .op(n10299) );
  nand2_1 U10537 ( .ip1(n11927), .ip2(\cache_data[11][25] ), .op(n10298) );
  nand2_1 U10538 ( .ip1(n11688), .ip2(\cache_data[14][25] ), .op(n10297) );
  nand4_1 U10539 ( .ip1(n10300), .ip2(n10299), .ip3(n10298), .ip4(n10297), 
        .op(n10317) );
  nand2_1 U10540 ( .ip1(n11966), .ip2(\cache_data[10][25] ), .op(n10304) );
  nand2_1 U10541 ( .ip1(n11964), .ip2(\cache_data[0][25] ), .op(n10303) );
  nand2_1 U10542 ( .ip1(n11943), .ip2(\cache_data[1][25] ), .op(n10302) );
  nand2_1 U10543 ( .ip1(n11973), .ip2(\cache_data[2][25] ), .op(n10301) );
  nand4_1 U10544 ( .ip1(n10304), .ip2(n10303), .ip3(n10302), .ip4(n10301), 
        .op(n10316) );
  nand2_1 U10545 ( .ip1(n12143), .ip2(\cache_data[7][25] ), .op(n10309) );
  nand2_1 U10546 ( .ip1(n12152), .ip2(\cache_data[9][25] ), .op(n10308) );
  nand2_1 U10547 ( .ip1(n10305), .ip2(\cache_data[6][25] ), .op(n10307) );
  nand2_1 U10548 ( .ip1(n12164), .ip2(\cache_data[4][25] ), .op(n10306) );
  nand4_1 U10549 ( .ip1(n10309), .ip2(n10308), .ip3(n10307), .ip4(n10306), 
        .op(n10315) );
  nand2_1 U10550 ( .ip1(n11965), .ip2(\cache_data[15][25] ), .op(n10313) );
  nand2_1 U10551 ( .ip1(n11963), .ip2(\cache_data[5][25] ), .op(n10312) );
  nand2_1 U10552 ( .ip1(n11978), .ip2(\cache_data[3][25] ), .op(n10311) );
  nand2_1 U10553 ( .ip1(n12191), .ip2(\cache_data[8][25] ), .op(n10310) );
  nand4_1 U10554 ( .ip1(n10313), .ip2(n10312), .ip3(n10311), .ip4(n10310), 
        .op(n10314) );
  or4_1 U10555 ( .ip1(n10317), .ip2(n10316), .ip3(n10315), .ip4(n10314), .op(
        n11243) );
  nand2_1 U10556 ( .ip1(n10828), .ip2(n11243), .op(n10382) );
  nand2_1 U10557 ( .ip1(n12164), .ip2(\cache_data[4][57] ), .op(n10321) );
  nand2_1 U10558 ( .ip1(n11963), .ip2(\cache_data[5][57] ), .op(n10320) );
  nand2_1 U10559 ( .ip1(n11927), .ip2(\cache_data[11][57] ), .op(n10319) );
  nand2_1 U10560 ( .ip1(n11964), .ip2(\cache_data[0][57] ), .op(n10318) );
  nand4_1 U10561 ( .ip1(n10321), .ip2(n10320), .ip3(n10319), .ip4(n10318), 
        .op(n10337) );
  nand2_1 U10562 ( .ip1(n12191), .ip2(\cache_data[8][57] ), .op(n10325) );
  nand2_1 U10563 ( .ip1(n11972), .ip2(\cache_data[6][57] ), .op(n10324) );
  nand2_1 U10564 ( .ip1(n12227), .ip2(\cache_data[12][57] ), .op(n10323) );
  nand2_1 U10565 ( .ip1(n11973), .ip2(\cache_data[2][57] ), .op(n10322) );
  nand4_1 U10566 ( .ip1(n10325), .ip2(n10324), .ip3(n10323), .ip4(n10322), 
        .op(n10336) );
  nand2_1 U10567 ( .ip1(n12165), .ip2(\cache_data[13][57] ), .op(n10329) );
  nand2_1 U10568 ( .ip1(n11978), .ip2(\cache_data[3][57] ), .op(n10328) );
  nand2_1 U10569 ( .ip1(n11943), .ip2(\cache_data[1][57] ), .op(n10327) );
  nand2_1 U10570 ( .ip1(n11688), .ip2(\cache_data[14][57] ), .op(n10326) );
  nand4_1 U10571 ( .ip1(n10329), .ip2(n10328), .ip3(n10327), .ip4(n10326), 
        .op(n10335) );
  nand2_1 U10572 ( .ip1(n11966), .ip2(\cache_data[10][57] ), .op(n10333) );
  nand2_1 U10573 ( .ip1(n12152), .ip2(\cache_data[9][57] ), .op(n10332) );
  nand2_1 U10574 ( .ip1(n11965), .ip2(\cache_data[15][57] ), .op(n10331) );
  nand2_1 U10575 ( .ip1(n12143), .ip2(\cache_data[7][57] ), .op(n10330) );
  nand4_1 U10576 ( .ip1(n10333), .ip2(n10332), .ip3(n10331), .ip4(n10330), 
        .op(n10334) );
  nor4_1 U10577 ( .ip1(n10337), .ip2(n10336), .ip3(n10335), .ip4(n10334), .op(
        n11240) );
  nor2_1 U10578 ( .ip1(n11240), .ip2(n10870), .op(n10359) );
  nand2_1 U10579 ( .ip1(n11963), .ip2(\cache_data[5][89] ), .op(n10341) );
  nand2_1 U10580 ( .ip1(n12152), .ip2(\cache_data[9][89] ), .op(n10340) );
  nand2_1 U10581 ( .ip1(n12143), .ip2(\cache_data[7][89] ), .op(n10339) );
  nand2_1 U10582 ( .ip1(n11966), .ip2(\cache_data[10][89] ), .op(n10338) );
  nand4_1 U10583 ( .ip1(n10341), .ip2(n10340), .ip3(n10339), .ip4(n10338), 
        .op(n10357) );
  nand2_1 U10584 ( .ip1(n11927), .ip2(\cache_data[11][89] ), .op(n10345) );
  nand2_1 U10585 ( .ip1(n11973), .ip2(\cache_data[2][89] ), .op(n10344) );
  nand2_1 U10586 ( .ip1(n11965), .ip2(\cache_data[15][89] ), .op(n10343) );
  nand2_1 U10587 ( .ip1(n12164), .ip2(\cache_data[4][89] ), .op(n10342) );
  nand4_1 U10588 ( .ip1(n10345), .ip2(n10344), .ip3(n10343), .ip4(n10342), 
        .op(n10356) );
  nand2_1 U10589 ( .ip1(n12165), .ip2(\cache_data[13][89] ), .op(n10349) );
  nand2_1 U10590 ( .ip1(n12227), .ip2(\cache_data[12][89] ), .op(n10348) );
  nand2_1 U10591 ( .ip1(n11972), .ip2(\cache_data[6][89] ), .op(n10347) );
  nand2_1 U10592 ( .ip1(n12191), .ip2(\cache_data[8][89] ), .op(n10346) );
  nand4_1 U10593 ( .ip1(n10349), .ip2(n10348), .ip3(n10347), .ip4(n10346), 
        .op(n10355) );
  nand2_1 U10594 ( .ip1(n11688), .ip2(\cache_data[14][89] ), .op(n10353) );
  nand2_1 U10595 ( .ip1(n11978), .ip2(\cache_data[3][89] ), .op(n10352) );
  nand2_1 U10596 ( .ip1(n11964), .ip2(\cache_data[0][89] ), .op(n10351) );
  nand2_1 U10597 ( .ip1(n11943), .ip2(\cache_data[1][89] ), .op(n10350) );
  nand4_1 U10598 ( .ip1(n10353), .ip2(n10352), .ip3(n10351), .ip4(n10350), 
        .op(n10354) );
  nor4_1 U10599 ( .ip1(n10357), .ip2(n10356), .ip3(n10355), .ip4(n10354), .op(
        n11239) );
  nor2_1 U10600 ( .ip1(n11239), .ip2(n10849), .op(n10358) );
  not_ab_or_c_or_d U10601 ( .ip1(data_wr_mem[25]), .ip2(n10873), .ip3(n10359), 
        .ip4(n10358), .op(n10381) );
  nand2_1 U10602 ( .ip1(n12164), .ip2(\cache_data[4][121] ), .op(n10363) );
  nand2_1 U10603 ( .ip1(n11688), .ip2(\cache_data[14][121] ), .op(n10362) );
  nand2_1 U10604 ( .ip1(n11965), .ip2(\cache_data[15][121] ), .op(n10361) );
  nand2_1 U10605 ( .ip1(n11963), .ip2(\cache_data[5][121] ), .op(n10360) );
  nand4_1 U10606 ( .ip1(n10363), .ip2(n10362), .ip3(n10361), .ip4(n10360), 
        .op(n10379) );
  nand2_1 U10607 ( .ip1(n11973), .ip2(\cache_data[2][121] ), .op(n10367) );
  nand2_1 U10608 ( .ip1(n11972), .ip2(\cache_data[6][121] ), .op(n10366) );
  nand2_1 U10609 ( .ip1(n11966), .ip2(\cache_data[10][121] ), .op(n10365) );
  nand2_1 U10610 ( .ip1(n12143), .ip2(\cache_data[7][121] ), .op(n10364) );
  nand4_1 U10611 ( .ip1(n10367), .ip2(n10366), .ip3(n10365), .ip4(n10364), 
        .op(n10378) );
  nand2_1 U10612 ( .ip1(n12191), .ip2(\cache_data[8][121] ), .op(n10371) );
  nand2_1 U10613 ( .ip1(n12227), .ip2(\cache_data[12][121] ), .op(n10370) );
  nand2_1 U10614 ( .ip1(n11943), .ip2(\cache_data[1][121] ), .op(n10369) );
  nand2_1 U10615 ( .ip1(n11927), .ip2(\cache_data[11][121] ), .op(n10368) );
  nand4_1 U10616 ( .ip1(n10371), .ip2(n10370), .ip3(n10369), .ip4(n10368), 
        .op(n10377) );
  nand2_1 U10617 ( .ip1(n12152), .ip2(\cache_data[9][121] ), .op(n10375) );
  nand2_1 U10618 ( .ip1(n11978), .ip2(\cache_data[3][121] ), .op(n10374) );
  nand2_1 U10619 ( .ip1(n11964), .ip2(\cache_data[0][121] ), .op(n10373) );
  nand2_1 U10620 ( .ip1(n12165), .ip2(\cache_data[13][121] ), .op(n10372) );
  nand4_1 U10621 ( .ip1(n10375), .ip2(n10374), .ip3(n10373), .ip4(n10372), 
        .op(n10376) );
  or4_1 U10622 ( .ip1(n10379), .ip2(n10378), .ip3(n10377), .ip4(n10376), .op(
        n11238) );
  nand2_1 U10623 ( .ip1(n10894), .ip2(n11238), .op(n10380) );
  nand3_1 U10624 ( .ip1(n10382), .ip2(n10381), .ip3(n10380), .op(n7423) );
  nand2_1 U10625 ( .ip1(n11966), .ip2(\cache_data[10][26] ), .op(n10386) );
  nand2_1 U10626 ( .ip1(n12152), .ip2(\cache_data[9][26] ), .op(n10385) );
  nand2_1 U10627 ( .ip1(n11972), .ip2(\cache_data[6][26] ), .op(n10384) );
  nand2_1 U10628 ( .ip1(n11973), .ip2(\cache_data[2][26] ), .op(n10383) );
  nand4_1 U10629 ( .ip1(n10386), .ip2(n10385), .ip3(n10384), .ip4(n10383), 
        .op(n10402) );
  nand2_1 U10630 ( .ip1(n12165), .ip2(\cache_data[13][26] ), .op(n10390) );
  nand2_1 U10631 ( .ip1(n12143), .ip2(\cache_data[7][26] ), .op(n10389) );
  nand2_1 U10632 ( .ip1(n11965), .ip2(\cache_data[15][26] ), .op(n10388) );
  nand2_1 U10633 ( .ip1(n11964), .ip2(\cache_data[0][26] ), .op(n10387) );
  nand4_1 U10634 ( .ip1(n10390), .ip2(n10389), .ip3(n10388), .ip4(n10387), 
        .op(n10401) );
  nand2_1 U10635 ( .ip1(n12164), .ip2(\cache_data[4][26] ), .op(n10394) );
  nand2_1 U10636 ( .ip1(n11943), .ip2(\cache_data[1][26] ), .op(n10393) );
  nand2_1 U10637 ( .ip1(n11978), .ip2(\cache_data[3][26] ), .op(n10392) );
  nand2_1 U10638 ( .ip1(n12191), .ip2(\cache_data[8][26] ), .op(n10391) );
  nand4_1 U10639 ( .ip1(n10394), .ip2(n10393), .ip3(n10392), .ip4(n10391), 
        .op(n10400) );
  nand2_1 U10640 ( .ip1(n11927), .ip2(\cache_data[11][26] ), .op(n10398) );
  nand2_1 U10641 ( .ip1(n12227), .ip2(\cache_data[12][26] ), .op(n10397) );
  nand2_1 U10642 ( .ip1(n11963), .ip2(\cache_data[5][26] ), .op(n10396) );
  nand2_1 U10643 ( .ip1(n11688), .ip2(\cache_data[14][26] ), .op(n10395) );
  nand4_1 U10644 ( .ip1(n10398), .ip2(n10397), .ip3(n10396), .ip4(n10395), 
        .op(n10399) );
  or4_1 U10645 ( .ip1(n10402), .ip2(n10401), .ip3(n10400), .ip4(n10399), .op(
        n11252) );
  nand2_1 U10646 ( .ip1(n10828), .ip2(n11252), .op(n10467) );
  nand2_1 U10647 ( .ip1(n11943), .ip2(\cache_data[1][90] ), .op(n10406) );
  nand2_1 U10648 ( .ip1(n11965), .ip2(\cache_data[15][90] ), .op(n10405) );
  nand2_1 U10649 ( .ip1(n12152), .ip2(\cache_data[9][90] ), .op(n10404) );
  nand2_1 U10650 ( .ip1(n12227), .ip2(\cache_data[12][90] ), .op(n10403) );
  nand4_1 U10651 ( .ip1(n10406), .ip2(n10405), .ip3(n10404), .ip4(n10403), 
        .op(n10422) );
  nand2_1 U10652 ( .ip1(n12165), .ip2(\cache_data[13][90] ), .op(n10410) );
  nand2_1 U10653 ( .ip1(n12164), .ip2(\cache_data[4][90] ), .op(n10409) );
  nand2_1 U10654 ( .ip1(n11966), .ip2(\cache_data[10][90] ), .op(n10408) );
  nand2_1 U10655 ( .ip1(n11927), .ip2(\cache_data[11][90] ), .op(n10407) );
  nand4_1 U10656 ( .ip1(n10410), .ip2(n10409), .ip3(n10408), .ip4(n10407), 
        .op(n10421) );
  nand2_1 U10657 ( .ip1(n11972), .ip2(\cache_data[6][90] ), .op(n10414) );
  nand2_1 U10658 ( .ip1(n11978), .ip2(\cache_data[3][90] ), .op(n10413) );
  nand2_1 U10659 ( .ip1(n11963), .ip2(\cache_data[5][90] ), .op(n10412) );
  nand2_1 U10660 ( .ip1(n11973), .ip2(\cache_data[2][90] ), .op(n10411) );
  nand4_1 U10661 ( .ip1(n10414), .ip2(n10413), .ip3(n10412), .ip4(n10411), 
        .op(n10420) );
  nand2_1 U10662 ( .ip1(n12143), .ip2(\cache_data[7][90] ), .op(n10418) );
  nand2_1 U10663 ( .ip1(n11964), .ip2(\cache_data[0][90] ), .op(n10417) );
  nand2_1 U10664 ( .ip1(n11688), .ip2(\cache_data[14][90] ), .op(n10416) );
  nand2_1 U10665 ( .ip1(n12191), .ip2(\cache_data[8][90] ), .op(n10415) );
  nand4_1 U10666 ( .ip1(n10418), .ip2(n10417), .ip3(n10416), .ip4(n10415), 
        .op(n10419) );
  nor4_1 U10667 ( .ip1(n10422), .ip2(n10421), .ip3(n10420), .ip4(n10419), .op(
        n11249) );
  nor2_1 U10668 ( .ip1(n11249), .ip2(n10849), .op(n10444) );
  nand2_1 U10669 ( .ip1(n12165), .ip2(\cache_data[13][58] ), .op(n10426) );
  nand2_1 U10670 ( .ip1(n12191), .ip2(\cache_data[8][58] ), .op(n10425) );
  nand2_1 U10671 ( .ip1(n11927), .ip2(\cache_data[11][58] ), .op(n10424) );
  nand2_1 U10672 ( .ip1(n11973), .ip2(\cache_data[2][58] ), .op(n10423) );
  nand4_1 U10673 ( .ip1(n10426), .ip2(n10425), .ip3(n10424), .ip4(n10423), 
        .op(n10442) );
  nand2_1 U10674 ( .ip1(n11978), .ip2(\cache_data[3][58] ), .op(n10430) );
  nand2_1 U10675 ( .ip1(n12143), .ip2(\cache_data[7][58] ), .op(n10429) );
  nand2_1 U10676 ( .ip1(n11688), .ip2(\cache_data[14][58] ), .op(n10428) );
  nand2_1 U10677 ( .ip1(n11972), .ip2(\cache_data[6][58] ), .op(n10427) );
  nand4_1 U10678 ( .ip1(n10430), .ip2(n10429), .ip3(n10428), .ip4(n10427), 
        .op(n10441) );
  nand2_1 U10679 ( .ip1(n11964), .ip2(\cache_data[0][58] ), .op(n10434) );
  nand2_1 U10680 ( .ip1(n12152), .ip2(\cache_data[9][58] ), .op(n10433) );
  nand2_1 U10681 ( .ip1(n11943), .ip2(\cache_data[1][58] ), .op(n10432) );
  nand2_1 U10682 ( .ip1(n11965), .ip2(\cache_data[15][58] ), .op(n10431) );
  nand4_1 U10683 ( .ip1(n10434), .ip2(n10433), .ip3(n10432), .ip4(n10431), 
        .op(n10440) );
  nand2_1 U10684 ( .ip1(n11966), .ip2(\cache_data[10][58] ), .op(n10438) );
  nand2_1 U10685 ( .ip1(n11963), .ip2(\cache_data[5][58] ), .op(n10437) );
  nand2_1 U10686 ( .ip1(n12227), .ip2(\cache_data[12][58] ), .op(n10436) );
  nand2_1 U10687 ( .ip1(n12164), .ip2(\cache_data[4][58] ), .op(n10435) );
  nand4_1 U10688 ( .ip1(n10438), .ip2(n10437), .ip3(n10436), .ip4(n10435), 
        .op(n10439) );
  nor4_1 U10689 ( .ip1(n10442), .ip2(n10441), .ip3(n10440), .ip4(n10439), .op(
        n11248) );
  nor2_1 U10690 ( .ip1(n11248), .ip2(n10870), .op(n10443) );
  not_ab_or_c_or_d U10691 ( .ip1(data_wr_mem[26]), .ip2(n10873), .ip3(n10444), 
        .ip4(n10443), .op(n10466) );
  nand2_1 U10692 ( .ip1(n12143), .ip2(\cache_data[7][122] ), .op(n10448) );
  nand2_1 U10693 ( .ip1(n12227), .ip2(\cache_data[12][122] ), .op(n10447) );
  nand2_1 U10694 ( .ip1(n12191), .ip2(\cache_data[8][122] ), .op(n10446) );
  nand2_1 U10695 ( .ip1(n11972), .ip2(\cache_data[6][122] ), .op(n10445) );
  nand4_1 U10696 ( .ip1(n10448), .ip2(n10447), .ip3(n10446), .ip4(n10445), 
        .op(n10464) );
  nand2_1 U10697 ( .ip1(n11978), .ip2(\cache_data[3][122] ), .op(n10452) );
  nand2_1 U10698 ( .ip1(n12152), .ip2(\cache_data[9][122] ), .op(n10451) );
  nand2_1 U10699 ( .ip1(n11964), .ip2(\cache_data[0][122] ), .op(n10450) );
  nand2_1 U10700 ( .ip1(n12164), .ip2(\cache_data[4][122] ), .op(n10449) );
  nand4_1 U10701 ( .ip1(n10452), .ip2(n10451), .ip3(n10450), .ip4(n10449), 
        .op(n10463) );
  nand2_1 U10702 ( .ip1(n11963), .ip2(\cache_data[5][122] ), .op(n10456) );
  nand2_1 U10703 ( .ip1(n11927), .ip2(\cache_data[11][122] ), .op(n10455) );
  nand2_1 U10704 ( .ip1(n11943), .ip2(\cache_data[1][122] ), .op(n10454) );
  nand2_1 U10705 ( .ip1(n11973), .ip2(\cache_data[2][122] ), .op(n10453) );
  nand4_1 U10706 ( .ip1(n10456), .ip2(n10455), .ip3(n10454), .ip4(n10453), 
        .op(n10462) );
  nand2_1 U10707 ( .ip1(n11688), .ip2(\cache_data[14][122] ), .op(n10460) );
  nand2_1 U10708 ( .ip1(n11965), .ip2(\cache_data[15][122] ), .op(n10459) );
  nand2_1 U10709 ( .ip1(n11966), .ip2(\cache_data[10][122] ), .op(n10458) );
  nand2_1 U10710 ( .ip1(n12165), .ip2(\cache_data[13][122] ), .op(n10457) );
  nand4_1 U10711 ( .ip1(n10460), .ip2(n10459), .ip3(n10458), .ip4(n10457), 
        .op(n10461) );
  or4_1 U10712 ( .ip1(n10464), .ip2(n10463), .ip3(n10462), .ip4(n10461), .op(
        n11247) );
  nand2_1 U10713 ( .ip1(n10894), .ip2(n11247), .op(n10465) );
  nand3_1 U10714 ( .ip1(n10467), .ip2(n10466), .ip3(n10465), .op(n7422) );
  nand2_1 U10715 ( .ip1(data_wr_mem[27]), .ip2(n10873), .op(n10552) );
  nand2_1 U10716 ( .ip1(n11972), .ip2(\cache_data[6][123] ), .op(n10471) );
  nand2_1 U10717 ( .ip1(n12242), .ip2(\cache_data[13][123] ), .op(n10470) );
  nand2_1 U10718 ( .ip1(n11964), .ip2(\cache_data[0][123] ), .op(n10469) );
  nand2_1 U10719 ( .ip1(n12234), .ip2(\cache_data[8][123] ), .op(n10468) );
  nand4_1 U10720 ( .ip1(n10471), .ip2(n10470), .ip3(n10469), .ip4(n10468), 
        .op(n10487) );
  nand2_1 U10721 ( .ip1(n11966), .ip2(\cache_data[10][123] ), .op(n10475) );
  nand2_1 U10722 ( .ip1(n11965), .ip2(\cache_data[15][123] ), .op(n10474) );
  nand2_1 U10723 ( .ip1(n11963), .ip2(\cache_data[5][123] ), .op(n10473) );
  nand2_1 U10724 ( .ip1(n12152), .ip2(\cache_data[9][123] ), .op(n10472) );
  nand4_1 U10725 ( .ip1(n10475), .ip2(n10474), .ip3(n10473), .ip4(n10472), 
        .op(n10486) );
  nand2_1 U10726 ( .ip1(n11973), .ip2(\cache_data[2][123] ), .op(n10479) );
  nand2_1 U10727 ( .ip1(n11688), .ip2(\cache_data[14][123] ), .op(n10478) );
  nand2_1 U10728 ( .ip1(n11978), .ip2(\cache_data[3][123] ), .op(n10477) );
  nand2_1 U10729 ( .ip1(n12170), .ip2(\cache_data[11][123] ), .op(n10476) );
  nand4_1 U10730 ( .ip1(n10479), .ip2(n10478), .ip3(n10477), .ip4(n10476), 
        .op(n10485) );
  nand2_1 U10731 ( .ip1(n12143), .ip2(\cache_data[7][123] ), .op(n10483) );
  nand2_1 U10732 ( .ip1(n12243), .ip2(\cache_data[4][123] ), .op(n10482) );
  inv_1 U10733 ( .ip(n11459), .op(n11979) );
  nand2_1 U10734 ( .ip1(n11979), .ip2(\cache_data[1][123] ), .op(n10481) );
  nand2_1 U10735 ( .ip1(n12030), .ip2(\cache_data[12][123] ), .op(n10480) );
  nand4_1 U10736 ( .ip1(n10483), .ip2(n10482), .ip3(n10481), .ip4(n10480), 
        .op(n10484) );
  or4_1 U10737 ( .ip1(n10487), .ip2(n10486), .ip3(n10485), .ip4(n10484), .op(
        n11256) );
  nand2_1 U10738 ( .ip1(n12242), .ip2(\cache_data[13][91] ), .op(n10491) );
  nand2_1 U10739 ( .ip1(n12152), .ip2(\cache_data[9][91] ), .op(n10490) );
  nand2_1 U10740 ( .ip1(n11978), .ip2(\cache_data[3][91] ), .op(n10489) );
  nand2_1 U10741 ( .ip1(n12243), .ip2(\cache_data[4][91] ), .op(n10488) );
  nand4_1 U10742 ( .ip1(n10491), .ip2(n10490), .ip3(n10489), .ip4(n10488), 
        .op(n10507) );
  nand2_1 U10743 ( .ip1(n12030), .ip2(\cache_data[12][91] ), .op(n10495) );
  nand2_1 U10744 ( .ip1(n11964), .ip2(\cache_data[0][91] ), .op(n10494) );
  nand2_1 U10745 ( .ip1(n11965), .ip2(\cache_data[15][91] ), .op(n10493) );
  nand2_1 U10746 ( .ip1(n11972), .ip2(\cache_data[6][91] ), .op(n10492) );
  nand4_1 U10747 ( .ip1(n10495), .ip2(n10494), .ip3(n10493), .ip4(n10492), 
        .op(n10506) );
  nand2_1 U10748 ( .ip1(n12234), .ip2(\cache_data[8][91] ), .op(n10499) );
  nand2_1 U10749 ( .ip1(n11688), .ip2(\cache_data[14][91] ), .op(n10498) );
  nand2_1 U10750 ( .ip1(n11973), .ip2(\cache_data[2][91] ), .op(n10497) );
  nand2_1 U10751 ( .ip1(n12143), .ip2(\cache_data[7][91] ), .op(n10496) );
  nand4_1 U10752 ( .ip1(n10499), .ip2(n10498), .ip3(n10497), .ip4(n10496), 
        .op(n10505) );
  nand2_1 U10753 ( .ip1(n11966), .ip2(\cache_data[10][91] ), .op(n10503) );
  nand2_1 U10754 ( .ip1(n12170), .ip2(\cache_data[11][91] ), .op(n10502) );
  nand2_1 U10755 ( .ip1(n11979), .ip2(\cache_data[1][91] ), .op(n10501) );
  nand2_1 U10756 ( .ip1(n11963), .ip2(\cache_data[5][91] ), .op(n10500) );
  nand4_1 U10757 ( .ip1(n10503), .ip2(n10502), .ip3(n10501), .ip4(n10500), 
        .op(n10504) );
  nor4_1 U10758 ( .ip1(n10507), .ip2(n10506), .ip3(n10505), .ip4(n10504), .op(
        n11258) );
  nor2_1 U10759 ( .ip1(n11258), .ip2(n10849), .op(n10529) );
  nand2_1 U10760 ( .ip1(n12234), .ip2(\cache_data[8][59] ), .op(n10511) );
  nand2_1 U10761 ( .ip1(n12243), .ip2(\cache_data[4][59] ), .op(n10510) );
  nand2_1 U10762 ( .ip1(n11966), .ip2(\cache_data[10][59] ), .op(n10509) );
  nand2_1 U10763 ( .ip1(n11978), .ip2(\cache_data[3][59] ), .op(n10508) );
  nand4_1 U10764 ( .ip1(n10511), .ip2(n10510), .ip3(n10509), .ip4(n10508), 
        .op(n10527) );
  nand2_1 U10765 ( .ip1(n12143), .ip2(\cache_data[7][59] ), .op(n10515) );
  nand2_1 U10766 ( .ip1(n11973), .ip2(\cache_data[2][59] ), .op(n10514) );
  nand2_1 U10767 ( .ip1(n11979), .ip2(\cache_data[1][59] ), .op(n10513) );
  nand2_1 U10768 ( .ip1(n12242), .ip2(\cache_data[13][59] ), .op(n10512) );
  nand4_1 U10769 ( .ip1(n10515), .ip2(n10514), .ip3(n10513), .ip4(n10512), 
        .op(n10526) );
  nand2_1 U10770 ( .ip1(n11972), .ip2(\cache_data[6][59] ), .op(n10519) );
  nand2_1 U10771 ( .ip1(n12030), .ip2(\cache_data[12][59] ), .op(n10518) );
  nand2_1 U10772 ( .ip1(n11963), .ip2(\cache_data[5][59] ), .op(n10517) );
  nand2_1 U10773 ( .ip1(n12170), .ip2(\cache_data[11][59] ), .op(n10516) );
  nand4_1 U10774 ( .ip1(n10519), .ip2(n10518), .ip3(n10517), .ip4(n10516), 
        .op(n10525) );
  nand2_1 U10775 ( .ip1(n11688), .ip2(\cache_data[14][59] ), .op(n10523) );
  nand2_1 U10776 ( .ip1(n11964), .ip2(\cache_data[0][59] ), .op(n10522) );
  nand2_1 U10777 ( .ip1(n11965), .ip2(\cache_data[15][59] ), .op(n10521) );
  nand2_1 U10778 ( .ip1(n12152), .ip2(\cache_data[9][59] ), .op(n10520) );
  nand4_1 U10779 ( .ip1(n10523), .ip2(n10522), .ip3(n10521), .ip4(n10520), 
        .op(n10524) );
  nor4_1 U10780 ( .ip1(n10527), .ip2(n10526), .ip3(n10525), .ip4(n10524), .op(
        n11257) );
  nor2_1 U10781 ( .ip1(n11257), .ip2(n10870), .op(n10528) );
  not_ab_or_c_or_d U10782 ( .ip1(n10894), .ip2(n11256), .ip3(n10529), .ip4(
        n10528), .op(n10551) );
  nand2_1 U10783 ( .ip1(n12170), .ip2(\cache_data[11][27] ), .op(n10533) );
  nand2_1 U10784 ( .ip1(n11979), .ip2(\cache_data[1][27] ), .op(n10532) );
  nand2_1 U10785 ( .ip1(n12242), .ip2(\cache_data[13][27] ), .op(n10531) );
  nand2_1 U10786 ( .ip1(n12152), .ip2(\cache_data[9][27] ), .op(n10530) );
  nand4_1 U10787 ( .ip1(n10533), .ip2(n10532), .ip3(n10531), .ip4(n10530), 
        .op(n10549) );
  nand2_1 U10788 ( .ip1(n12234), .ip2(\cache_data[8][27] ), .op(n10537) );
  nand2_1 U10789 ( .ip1(n11972), .ip2(\cache_data[6][27] ), .op(n10536) );
  nand2_1 U10790 ( .ip1(n12030), .ip2(\cache_data[12][27] ), .op(n10535) );
  nand2_1 U10791 ( .ip1(n11966), .ip2(\cache_data[10][27] ), .op(n10534) );
  nand4_1 U10792 ( .ip1(n10537), .ip2(n10536), .ip3(n10535), .ip4(n10534), 
        .op(n10548) );
  nand2_1 U10793 ( .ip1(n11963), .ip2(\cache_data[5][27] ), .op(n10541) );
  nand2_1 U10794 ( .ip1(n11965), .ip2(\cache_data[15][27] ), .op(n10540) );
  nand2_1 U10795 ( .ip1(n11688), .ip2(\cache_data[14][27] ), .op(n10539) );
  nand2_1 U10796 ( .ip1(n11973), .ip2(\cache_data[2][27] ), .op(n10538) );
  nand4_1 U10797 ( .ip1(n10541), .ip2(n10540), .ip3(n10539), .ip4(n10538), 
        .op(n10547) );
  nand2_1 U10798 ( .ip1(n12243), .ip2(\cache_data[4][27] ), .op(n10545) );
  nand2_1 U10799 ( .ip1(n11978), .ip2(\cache_data[3][27] ), .op(n10544) );
  nand2_1 U10800 ( .ip1(n12143), .ip2(\cache_data[7][27] ), .op(n10543) );
  nand2_1 U10801 ( .ip1(n11964), .ip2(\cache_data[0][27] ), .op(n10542) );
  nand4_1 U10802 ( .ip1(n10545), .ip2(n10544), .ip3(n10543), .ip4(n10542), 
        .op(n10546) );
  or4_1 U10803 ( .ip1(n10549), .ip2(n10548), .ip3(n10547), .ip4(n10546), .op(
        n11261) );
  nand2_1 U10804 ( .ip1(n10828), .ip2(n11261), .op(n10550) );
  nand3_1 U10805 ( .ip1(n10552), .ip2(n10551), .ip3(n10550), .op(n7421) );
  nand2_1 U10806 ( .ip1(n12242), .ip2(\cache_data[13][28] ), .op(n10556) );
  nand2_1 U10807 ( .ip1(n11979), .ip2(\cache_data[1][28] ), .op(n10555) );
  nand2_1 U10808 ( .ip1(n12170), .ip2(\cache_data[11][28] ), .op(n10554) );
  nand2_1 U10809 ( .ip1(n11688), .ip2(\cache_data[14][28] ), .op(n10553) );
  nand4_1 U10810 ( .ip1(n10556), .ip2(n10555), .ip3(n10554), .ip4(n10553), 
        .op(n10572) );
  nand2_1 U10811 ( .ip1(n11964), .ip2(\cache_data[0][28] ), .op(n10560) );
  nand2_1 U10812 ( .ip1(n11978), .ip2(\cache_data[3][28] ), .op(n10559) );
  nand2_1 U10813 ( .ip1(n11963), .ip2(\cache_data[5][28] ), .op(n10558) );
  nand2_1 U10814 ( .ip1(n12152), .ip2(\cache_data[9][28] ), .op(n10557) );
  nand4_1 U10815 ( .ip1(n10560), .ip2(n10559), .ip3(n10558), .ip4(n10557), 
        .op(n10571) );
  nand2_1 U10816 ( .ip1(n11965), .ip2(\cache_data[15][28] ), .op(n10564) );
  nand2_1 U10817 ( .ip1(n12234), .ip2(\cache_data[8][28] ), .op(n10563) );
  nand2_1 U10818 ( .ip1(n11973), .ip2(\cache_data[2][28] ), .op(n10562) );
  nand2_1 U10819 ( .ip1(n12143), .ip2(\cache_data[7][28] ), .op(n10561) );
  nand4_1 U10820 ( .ip1(n10564), .ip2(n10563), .ip3(n10562), .ip4(n10561), 
        .op(n10570) );
  nand2_1 U10821 ( .ip1(n11966), .ip2(\cache_data[10][28] ), .op(n10568) );
  nand2_1 U10822 ( .ip1(n11972), .ip2(\cache_data[6][28] ), .op(n10567) );
  nand2_1 U10823 ( .ip1(n12243), .ip2(\cache_data[4][28] ), .op(n10566) );
  nand2_1 U10824 ( .ip1(n12030), .ip2(\cache_data[12][28] ), .op(n10565) );
  nand4_1 U10825 ( .ip1(n10568), .ip2(n10567), .ip3(n10566), .ip4(n10565), 
        .op(n10569) );
  or4_1 U10826 ( .ip1(n10572), .ip2(n10571), .ip3(n10570), .ip4(n10569), .op(
        n11270) );
  nand2_1 U10827 ( .ip1(n10828), .ip2(n11270), .op(n10637) );
  nand2_1 U10828 ( .ip1(n11978), .ip2(\cache_data[3][92] ), .op(n10576) );
  nand2_1 U10829 ( .ip1(n12170), .ip2(\cache_data[11][92] ), .op(n10575) );
  nand2_1 U10830 ( .ip1(n11973), .ip2(\cache_data[2][92] ), .op(n10574) );
  nand2_1 U10831 ( .ip1(n12152), .ip2(\cache_data[9][92] ), .op(n10573) );
  nand4_1 U10832 ( .ip1(n10576), .ip2(n10575), .ip3(n10574), .ip4(n10573), 
        .op(n10592) );
  nand2_1 U10833 ( .ip1(n11963), .ip2(\cache_data[5][92] ), .op(n10580) );
  nand2_1 U10834 ( .ip1(n11688), .ip2(\cache_data[14][92] ), .op(n10579) );
  nand2_1 U10835 ( .ip1(n12243), .ip2(\cache_data[4][92] ), .op(n10578) );
  nand2_1 U10836 ( .ip1(n12234), .ip2(\cache_data[8][92] ), .op(n10577) );
  nand4_1 U10837 ( .ip1(n10580), .ip2(n10579), .ip3(n10578), .ip4(n10577), 
        .op(n10591) );
  nand2_1 U10838 ( .ip1(n11972), .ip2(\cache_data[6][92] ), .op(n10584) );
  nand2_1 U10839 ( .ip1(n11966), .ip2(\cache_data[10][92] ), .op(n10583) );
  nand2_1 U10840 ( .ip1(n11965), .ip2(\cache_data[15][92] ), .op(n10582) );
  nand2_1 U10841 ( .ip1(n12030), .ip2(\cache_data[12][92] ), .op(n10581) );
  nand4_1 U10842 ( .ip1(n10584), .ip2(n10583), .ip3(n10582), .ip4(n10581), 
        .op(n10590) );
  nand2_1 U10843 ( .ip1(n11964), .ip2(\cache_data[0][92] ), .op(n10588) );
  nand2_1 U10844 ( .ip1(n12242), .ip2(\cache_data[13][92] ), .op(n10587) );
  nand2_1 U10845 ( .ip1(n11979), .ip2(\cache_data[1][92] ), .op(n10586) );
  nand2_1 U10846 ( .ip1(n12143), .ip2(\cache_data[7][92] ), .op(n10585) );
  nand4_1 U10847 ( .ip1(n10588), .ip2(n10587), .ip3(n10586), .ip4(n10585), 
        .op(n10589) );
  nor4_1 U10848 ( .ip1(n10592), .ip2(n10591), .ip3(n10590), .ip4(n10589), .op(
        n11267) );
  nor2_1 U10849 ( .ip1(n11267), .ip2(n10849), .op(n10614) );
  nand2_1 U10850 ( .ip1(n11963), .ip2(\cache_data[5][60] ), .op(n10596) );
  nand2_1 U10851 ( .ip1(n11972), .ip2(\cache_data[6][60] ), .op(n10595) );
  nand2_1 U10852 ( .ip1(n11964), .ip2(\cache_data[0][60] ), .op(n10594) );
  nand2_1 U10853 ( .ip1(n11966), .ip2(\cache_data[10][60] ), .op(n10593) );
  nand4_1 U10854 ( .ip1(n10596), .ip2(n10595), .ip3(n10594), .ip4(n10593), 
        .op(n10612) );
  nand2_1 U10855 ( .ip1(n12243), .ip2(\cache_data[4][60] ), .op(n10600) );
  nand2_1 U10856 ( .ip1(n11688), .ip2(\cache_data[14][60] ), .op(n10599) );
  nand2_1 U10857 ( .ip1(n12242), .ip2(\cache_data[13][60] ), .op(n10598) );
  nand2_1 U10858 ( .ip1(n12143), .ip2(\cache_data[7][60] ), .op(n10597) );
  nand4_1 U10859 ( .ip1(n10600), .ip2(n10599), .ip3(n10598), .ip4(n10597), 
        .op(n10611) );
  nand2_1 U10860 ( .ip1(n12170), .ip2(\cache_data[11][60] ), .op(n10604) );
  nand2_1 U10861 ( .ip1(n11965), .ip2(\cache_data[15][60] ), .op(n10603) );
  nand2_1 U10862 ( .ip1(n12152), .ip2(\cache_data[9][60] ), .op(n10602) );
  nand2_1 U10863 ( .ip1(n11973), .ip2(\cache_data[2][60] ), .op(n10601) );
  nand4_1 U10864 ( .ip1(n10604), .ip2(n10603), .ip3(n10602), .ip4(n10601), 
        .op(n10610) );
  nand2_1 U10865 ( .ip1(n11978), .ip2(\cache_data[3][60] ), .op(n10608) );
  nand2_1 U10866 ( .ip1(n12234), .ip2(\cache_data[8][60] ), .op(n10607) );
  nand2_1 U10867 ( .ip1(n11979), .ip2(\cache_data[1][60] ), .op(n10606) );
  nand2_1 U10868 ( .ip1(n12030), .ip2(\cache_data[12][60] ), .op(n10605) );
  nand4_1 U10869 ( .ip1(n10608), .ip2(n10607), .ip3(n10606), .ip4(n10605), 
        .op(n10609) );
  nor4_1 U10870 ( .ip1(n10612), .ip2(n10611), .ip3(n10610), .ip4(n10609), .op(
        n11266) );
  nor2_1 U10871 ( .ip1(n11266), .ip2(n10870), .op(n10613) );
  not_ab_or_c_or_d U10872 ( .ip1(data_wr_mem[28]), .ip2(n10873), .ip3(n10614), 
        .ip4(n10613), .op(n10636) );
  nand2_1 U10873 ( .ip1(n11964), .ip2(\cache_data[0][124] ), .op(n10618) );
  nand2_1 U10874 ( .ip1(n11973), .ip2(\cache_data[2][124] ), .op(n10617) );
  nand2_1 U10875 ( .ip1(n11978), .ip2(\cache_data[3][124] ), .op(n10616) );
  nand2_1 U10876 ( .ip1(n11963), .ip2(\cache_data[5][124] ), .op(n10615) );
  nand4_1 U10877 ( .ip1(n10618), .ip2(n10617), .ip3(n10616), .ip4(n10615), 
        .op(n10634) );
  nand2_1 U10878 ( .ip1(n11972), .ip2(\cache_data[6][124] ), .op(n10622) );
  nand2_1 U10879 ( .ip1(n12152), .ip2(\cache_data[9][124] ), .op(n10621) );
  nand2_1 U10880 ( .ip1(n12143), .ip2(\cache_data[7][124] ), .op(n10620) );
  nand2_1 U10881 ( .ip1(n12030), .ip2(\cache_data[12][124] ), .op(n10619) );
  nand4_1 U10882 ( .ip1(n10622), .ip2(n10621), .ip3(n10620), .ip4(n10619), 
        .op(n10633) );
  nand2_1 U10883 ( .ip1(n11979), .ip2(\cache_data[1][124] ), .op(n10626) );
  nand2_1 U10884 ( .ip1(n11966), .ip2(\cache_data[10][124] ), .op(n10625) );
  nand2_1 U10885 ( .ip1(n12170), .ip2(\cache_data[11][124] ), .op(n10624) );
  nand2_1 U10886 ( .ip1(n11965), .ip2(\cache_data[15][124] ), .op(n10623) );
  nand4_1 U10887 ( .ip1(n10626), .ip2(n10625), .ip3(n10624), .ip4(n10623), 
        .op(n10632) );
  nand2_1 U10888 ( .ip1(n12234), .ip2(\cache_data[8][124] ), .op(n10630) );
  nand2_1 U10889 ( .ip1(n12243), .ip2(\cache_data[4][124] ), .op(n10629) );
  nand2_1 U10890 ( .ip1(n11688), .ip2(\cache_data[14][124] ), .op(n10628) );
  nand2_1 U10891 ( .ip1(n12242), .ip2(\cache_data[13][124] ), .op(n10627) );
  nand4_1 U10892 ( .ip1(n10630), .ip2(n10629), .ip3(n10628), .ip4(n10627), 
        .op(n10631) );
  or4_1 U10893 ( .ip1(n10634), .ip2(n10633), .ip3(n10632), .ip4(n10631), .op(
        n11265) );
  nand2_1 U10894 ( .ip1(n10894), .ip2(n11265), .op(n10635) );
  nand3_1 U10895 ( .ip1(n10637), .ip2(n10636), .ip3(n10635), .op(n7420) );
  nand2_1 U10896 ( .ip1(n12243), .ip2(\cache_data[4][29] ), .op(n10641) );
  nand2_1 U10897 ( .ip1(n11965), .ip2(\cache_data[15][29] ), .op(n10640) );
  nand2_1 U10898 ( .ip1(n11973), .ip2(\cache_data[2][29] ), .op(n10639) );
  nand2_1 U10899 ( .ip1(n12242), .ip2(\cache_data[13][29] ), .op(n10638) );
  nand4_1 U10900 ( .ip1(n10641), .ip2(n10640), .ip3(n10639), .ip4(n10638), 
        .op(n10657) );
  nand2_1 U10901 ( .ip1(n12170), .ip2(\cache_data[11][29] ), .op(n10645) );
  nand2_1 U10902 ( .ip1(n11964), .ip2(\cache_data[0][29] ), .op(n10644) );
  nand2_1 U10903 ( .ip1(n11688), .ip2(\cache_data[14][29] ), .op(n10643) );
  nand2_1 U10904 ( .ip1(n11963), .ip2(\cache_data[5][29] ), .op(n10642) );
  nand4_1 U10905 ( .ip1(n10645), .ip2(n10644), .ip3(n10643), .ip4(n10642), 
        .op(n10656) );
  nand2_1 U10906 ( .ip1(n11972), .ip2(\cache_data[6][29] ), .op(n10649) );
  nand2_1 U10907 ( .ip1(n12030), .ip2(\cache_data[12][29] ), .op(n10648) );
  nand2_1 U10908 ( .ip1(n11979), .ip2(\cache_data[1][29] ), .op(n10647) );
  nand2_1 U10909 ( .ip1(n12234), .ip2(\cache_data[8][29] ), .op(n10646) );
  nand4_1 U10910 ( .ip1(n10649), .ip2(n10648), .ip3(n10647), .ip4(n10646), 
        .op(n10655) );
  nand2_1 U10911 ( .ip1(n11966), .ip2(\cache_data[10][29] ), .op(n10653) );
  nand2_1 U10912 ( .ip1(n12152), .ip2(\cache_data[9][29] ), .op(n10652) );
  nand2_1 U10913 ( .ip1(n11978), .ip2(\cache_data[3][29] ), .op(n10651) );
  nand2_1 U10914 ( .ip1(n12143), .ip2(\cache_data[7][29] ), .op(n10650) );
  nand4_1 U10915 ( .ip1(n10653), .ip2(n10652), .ip3(n10651), .ip4(n10650), 
        .op(n10654) );
  or4_1 U10916 ( .ip1(n10657), .ip2(n10656), .ip3(n10655), .ip4(n10654), .op(
        n11279) );
  nand2_1 U10917 ( .ip1(n10828), .ip2(n11279), .op(n10722) );
  nand2_1 U10918 ( .ip1(n11973), .ip2(\cache_data[2][61] ), .op(n10661) );
  nand2_1 U10919 ( .ip1(n11979), .ip2(\cache_data[1][61] ), .op(n10660) );
  nand2_1 U10920 ( .ip1(n11978), .ip2(\cache_data[3][61] ), .op(n10659) );
  nand2_1 U10921 ( .ip1(n12242), .ip2(\cache_data[13][61] ), .op(n10658) );
  nand4_1 U10922 ( .ip1(n10661), .ip2(n10660), .ip3(n10659), .ip4(n10658), 
        .op(n10677) );
  nand2_1 U10923 ( .ip1(n12152), .ip2(\cache_data[9][61] ), .op(n10665) );
  nand2_1 U10924 ( .ip1(n11964), .ip2(\cache_data[0][61] ), .op(n10664) );
  nand2_1 U10925 ( .ip1(n12143), .ip2(\cache_data[7][61] ), .op(n10663) );
  nand2_1 U10926 ( .ip1(n12234), .ip2(\cache_data[8][61] ), .op(n10662) );
  nand4_1 U10927 ( .ip1(n10665), .ip2(n10664), .ip3(n10663), .ip4(n10662), 
        .op(n10676) );
  nand2_1 U10928 ( .ip1(n11972), .ip2(\cache_data[6][61] ), .op(n10669) );
  nand2_1 U10929 ( .ip1(n11966), .ip2(\cache_data[10][61] ), .op(n10668) );
  nand2_1 U10930 ( .ip1(n12030), .ip2(\cache_data[12][61] ), .op(n10667) );
  nand2_1 U10931 ( .ip1(n12170), .ip2(\cache_data[11][61] ), .op(n10666) );
  nand4_1 U10932 ( .ip1(n10669), .ip2(n10668), .ip3(n10667), .ip4(n10666), 
        .op(n10675) );
  nand2_1 U10933 ( .ip1(n12243), .ip2(\cache_data[4][61] ), .op(n10673) );
  nand2_1 U10934 ( .ip1(n11963), .ip2(\cache_data[5][61] ), .op(n10672) );
  nand2_1 U10935 ( .ip1(n11688), .ip2(\cache_data[14][61] ), .op(n10671) );
  nand2_1 U10936 ( .ip1(n11965), .ip2(\cache_data[15][61] ), .op(n10670) );
  nand4_1 U10937 ( .ip1(n10673), .ip2(n10672), .ip3(n10671), .ip4(n10670), 
        .op(n10674) );
  nor4_1 U10938 ( .ip1(n10677), .ip2(n10676), .ip3(n10675), .ip4(n10674), .op(
        n11275) );
  nor2_1 U10939 ( .ip1(n11275), .ip2(n10870), .op(n10699) );
  nand2_1 U10940 ( .ip1(n11978), .ip2(\cache_data[3][93] ), .op(n10681) );
  nand2_1 U10941 ( .ip1(n11979), .ip2(\cache_data[1][93] ), .op(n10680) );
  nand2_1 U10942 ( .ip1(n11973), .ip2(\cache_data[2][93] ), .op(n10679) );
  nand2_1 U10943 ( .ip1(n11688), .ip2(\cache_data[14][93] ), .op(n10678) );
  nand4_1 U10944 ( .ip1(n10681), .ip2(n10680), .ip3(n10679), .ip4(n10678), 
        .op(n10697) );
  nand2_1 U10945 ( .ip1(n11964), .ip2(\cache_data[0][93] ), .op(n10685) );
  nand2_1 U10946 ( .ip1(n12170), .ip2(\cache_data[11][93] ), .op(n10684) );
  nand2_1 U10947 ( .ip1(n11972), .ip2(\cache_data[6][93] ), .op(n10683) );
  nand2_1 U10948 ( .ip1(n12030), .ip2(\cache_data[12][93] ), .op(n10682) );
  nand4_1 U10949 ( .ip1(n10685), .ip2(n10684), .ip3(n10683), .ip4(n10682), 
        .op(n10696) );
  nand2_1 U10950 ( .ip1(n11963), .ip2(\cache_data[5][93] ), .op(n10689) );
  nand2_1 U10951 ( .ip1(n12143), .ip2(\cache_data[7][93] ), .op(n10688) );
  nand2_1 U10952 ( .ip1(n12152), .ip2(\cache_data[9][93] ), .op(n10687) );
  nand2_1 U10953 ( .ip1(n11965), .ip2(\cache_data[15][93] ), .op(n10686) );
  nand4_1 U10954 ( .ip1(n10689), .ip2(n10688), .ip3(n10687), .ip4(n10686), 
        .op(n10695) );
  nand2_1 U10955 ( .ip1(n12242), .ip2(\cache_data[13][93] ), .op(n10693) );
  nand2_1 U10956 ( .ip1(n11966), .ip2(\cache_data[10][93] ), .op(n10692) );
  nand2_1 U10957 ( .ip1(n12234), .ip2(\cache_data[8][93] ), .op(n10691) );
  nand2_1 U10958 ( .ip1(n12243), .ip2(\cache_data[4][93] ), .op(n10690) );
  nand4_1 U10959 ( .ip1(n10693), .ip2(n10692), .ip3(n10691), .ip4(n10690), 
        .op(n10694) );
  nor4_1 U10960 ( .ip1(n10697), .ip2(n10696), .ip3(n10695), .ip4(n10694), .op(
        n11276) );
  nor2_1 U10961 ( .ip1(n11276), .ip2(n10849), .op(n10698) );
  not_ab_or_c_or_d U10962 ( .ip1(data_wr_mem[29]), .ip2(n10873), .ip3(n10699), 
        .ip4(n10698), .op(n10721) );
  nand2_1 U10963 ( .ip1(n12143), .ip2(\cache_data[7][125] ), .op(n10703) );
  nand2_1 U10964 ( .ip1(n11688), .ip2(\cache_data[14][125] ), .op(n10702) );
  nand2_1 U10965 ( .ip1(n12170), .ip2(\cache_data[11][125] ), .op(n10701) );
  nand2_1 U10966 ( .ip1(n11972), .ip2(\cache_data[6][125] ), .op(n10700) );
  nand4_1 U10967 ( .ip1(n10703), .ip2(n10702), .ip3(n10701), .ip4(n10700), 
        .op(n10719) );
  nand2_1 U10968 ( .ip1(n11978), .ip2(\cache_data[3][125] ), .op(n10707) );
  nand2_1 U10969 ( .ip1(n12243), .ip2(\cache_data[4][125] ), .op(n10706) );
  nand2_1 U10970 ( .ip1(n11963), .ip2(\cache_data[5][125] ), .op(n10705) );
  nand2_1 U10971 ( .ip1(n11966), .ip2(\cache_data[10][125] ), .op(n10704) );
  nand4_1 U10972 ( .ip1(n10707), .ip2(n10706), .ip3(n10705), .ip4(n10704), 
        .op(n10718) );
  nand2_1 U10973 ( .ip1(n11965), .ip2(\cache_data[15][125] ), .op(n10711) );
  nand2_1 U10974 ( .ip1(n12234), .ip2(\cache_data[8][125] ), .op(n10710) );
  nand2_1 U10975 ( .ip1(n12152), .ip2(\cache_data[9][125] ), .op(n10709) );
  nand2_1 U10976 ( .ip1(n11964), .ip2(\cache_data[0][125] ), .op(n10708) );
  nand4_1 U10977 ( .ip1(n10711), .ip2(n10710), .ip3(n10709), .ip4(n10708), 
        .op(n10717) );
  nand2_1 U10978 ( .ip1(n11973), .ip2(\cache_data[2][125] ), .op(n10715) );
  nand2_1 U10979 ( .ip1(n12030), .ip2(\cache_data[12][125] ), .op(n10714) );
  nand2_1 U10980 ( .ip1(n11979), .ip2(\cache_data[1][125] ), .op(n10713) );
  nand2_1 U10981 ( .ip1(n12242), .ip2(\cache_data[13][125] ), .op(n10712) );
  nand4_1 U10982 ( .ip1(n10715), .ip2(n10714), .ip3(n10713), .ip4(n10712), 
        .op(n10716) );
  or4_1 U10983 ( .ip1(n10719), .ip2(n10718), .ip3(n10717), .ip4(n10716), .op(
        n11274) );
  nand2_1 U10984 ( .ip1(n10894), .ip2(n11274), .op(n10720) );
  nand3_1 U10985 ( .ip1(n10722), .ip2(n10721), .ip3(n10720), .op(n7419) );
  nand2_1 U10986 ( .ip1(data_wr_mem[30]), .ip2(n10873), .op(n10807) );
  nand2_1 U10987 ( .ip1(n12241), .ip2(\cache_data[9][30] ), .op(n10726) );
  nand2_1 U10988 ( .ip1(n11979), .ip2(\cache_data[1][30] ), .op(n10725) );
  nand2_1 U10989 ( .ip1(n11965), .ip2(\cache_data[15][30] ), .op(n10724) );
  nand2_1 U10990 ( .ip1(n12242), .ip2(\cache_data[13][30] ), .op(n10723) );
  nand4_1 U10991 ( .ip1(n10726), .ip2(n10725), .ip3(n10724), .ip4(n10723), 
        .op(n10742) );
  nand2_1 U10992 ( .ip1(n12202), .ip2(\cache_data[7][30] ), .op(n10730) );
  nand2_1 U10993 ( .ip1(n11964), .ip2(\cache_data[0][30] ), .op(n10729) );
  nand2_1 U10994 ( .ip1(n12164), .ip2(\cache_data[4][30] ), .op(n10728) );
  nand2_1 U10995 ( .ip1(n11972), .ip2(\cache_data[6][30] ), .op(n10727) );
  nand4_1 U10996 ( .ip1(n10730), .ip2(n10729), .ip3(n10728), .ip4(n10727), 
        .op(n10741) );
  nand2_1 U10997 ( .ip1(n11688), .ip2(\cache_data[14][30] ), .op(n10734) );
  nand2_1 U10998 ( .ip1(n11963), .ip2(\cache_data[5][30] ), .op(n10733) );
  nand2_1 U10999 ( .ip1(n11978), .ip2(\cache_data[3][30] ), .op(n10732) );
  nand2_1 U11000 ( .ip1(n12170), .ip2(\cache_data[11][30] ), .op(n10731) );
  nand4_1 U11001 ( .ip1(n10734), .ip2(n10733), .ip3(n10732), .ip4(n10731), 
        .op(n10740) );
  nand2_1 U11002 ( .ip1(n11973), .ip2(\cache_data[2][30] ), .op(n10738) );
  nand2_1 U11003 ( .ip1(n12234), .ip2(\cache_data[8][30] ), .op(n10737) );
  nand2_1 U11004 ( .ip1(n12030), .ip2(\cache_data[12][30] ), .op(n10736) );
  nand2_1 U11005 ( .ip1(n11966), .ip2(\cache_data[10][30] ), .op(n10735) );
  nand4_1 U11006 ( .ip1(n10738), .ip2(n10737), .ip3(n10736), .ip4(n10735), 
        .op(n10739) );
  or4_1 U11007 ( .ip1(n10742), .ip2(n10741), .ip3(n10740), .ip4(n10739), .op(
        n11283) );
  nand2_1 U11008 ( .ip1(n12202), .ip2(\cache_data[7][94] ), .op(n10746) );
  nand2_1 U11009 ( .ip1(n12170), .ip2(\cache_data[11][94] ), .op(n10745) );
  nand2_1 U11010 ( .ip1(n11964), .ip2(\cache_data[0][94] ), .op(n10744) );
  nand2_1 U11011 ( .ip1(n11943), .ip2(\cache_data[1][94] ), .op(n10743) );
  nand4_1 U11012 ( .ip1(n10746), .ip2(n10745), .ip3(n10744), .ip4(n10743), 
        .op(n10762) );
  nand2_1 U11013 ( .ip1(n12164), .ip2(\cache_data[4][94] ), .op(n10750) );
  nand2_1 U11014 ( .ip1(n11973), .ip2(\cache_data[2][94] ), .op(n10749) );
  nand2_1 U11015 ( .ip1(n11966), .ip2(\cache_data[10][94] ), .op(n10748) );
  nand2_1 U11016 ( .ip1(n12242), .ip2(\cache_data[13][94] ), .op(n10747) );
  nand4_1 U11017 ( .ip1(n10750), .ip2(n10749), .ip3(n10748), .ip4(n10747), 
        .op(n10761) );
  nand2_1 U11018 ( .ip1(n11978), .ip2(\cache_data[3][94] ), .op(n10754) );
  nand2_1 U11019 ( .ip1(n11963), .ip2(\cache_data[5][94] ), .op(n10753) );
  nand2_1 U11020 ( .ip1(n12234), .ip2(\cache_data[8][94] ), .op(n10752) );
  nand2_1 U11021 ( .ip1(n12241), .ip2(\cache_data[9][94] ), .op(n10751) );
  nand4_1 U11022 ( .ip1(n10754), .ip2(n10753), .ip3(n10752), .ip4(n10751), 
        .op(n10760) );
  nand2_1 U11023 ( .ip1(n11965), .ip2(\cache_data[15][94] ), .op(n10758) );
  nand2_1 U11024 ( .ip1(n11972), .ip2(\cache_data[6][94] ), .op(n10757) );
  nand2_1 U11025 ( .ip1(n12030), .ip2(\cache_data[12][94] ), .op(n10756) );
  nand2_1 U11026 ( .ip1(n11688), .ip2(\cache_data[14][94] ), .op(n10755) );
  nand4_1 U11027 ( .ip1(n10758), .ip2(n10757), .ip3(n10756), .ip4(n10755), 
        .op(n10759) );
  nor4_1 U11028 ( .ip1(n10762), .ip2(n10761), .ip3(n10760), .ip4(n10759), .op(
        n11285) );
  nor2_1 U11029 ( .ip1(n11285), .ip2(n10849), .op(n10784) );
  nand2_1 U11030 ( .ip1(n11966), .ip2(\cache_data[10][62] ), .op(n10766) );
  nand2_1 U11031 ( .ip1(n12202), .ip2(\cache_data[7][62] ), .op(n10765) );
  nand2_1 U11032 ( .ip1(n12170), .ip2(\cache_data[11][62] ), .op(n10764) );
  nand2_1 U11033 ( .ip1(n11972), .ip2(\cache_data[6][62] ), .op(n10763) );
  nand4_1 U11034 ( .ip1(n10766), .ip2(n10765), .ip3(n10764), .ip4(n10763), 
        .op(n10782) );
  nand2_1 U11035 ( .ip1(n11973), .ip2(\cache_data[2][62] ), .op(n10770) );
  nand2_1 U11036 ( .ip1(n12242), .ip2(\cache_data[13][62] ), .op(n10769) );
  nand2_1 U11037 ( .ip1(n11963), .ip2(\cache_data[5][62] ), .op(n10768) );
  nand2_1 U11038 ( .ip1(n11964), .ip2(\cache_data[0][62] ), .op(n10767) );
  nand4_1 U11039 ( .ip1(n10770), .ip2(n10769), .ip3(n10768), .ip4(n10767), 
        .op(n10781) );
  nand2_1 U11040 ( .ip1(n11965), .ip2(\cache_data[15][62] ), .op(n10774) );
  nand2_1 U11041 ( .ip1(n12241), .ip2(\cache_data[9][62] ), .op(n10773) );
  nand2_1 U11042 ( .ip1(n11978), .ip2(\cache_data[3][62] ), .op(n10772) );
  nand2_1 U11043 ( .ip1(n12234), .ip2(\cache_data[8][62] ), .op(n10771) );
  nand4_1 U11044 ( .ip1(n10774), .ip2(n10773), .ip3(n10772), .ip4(n10771), 
        .op(n10780) );
  nand2_1 U11045 ( .ip1(n11979), .ip2(\cache_data[1][62] ), .op(n10778) );
  nand2_1 U11046 ( .ip1(n11688), .ip2(\cache_data[14][62] ), .op(n10777) );
  nand2_1 U11047 ( .ip1(n12030), .ip2(\cache_data[12][62] ), .op(n10776) );
  nand2_1 U11048 ( .ip1(n12164), .ip2(\cache_data[4][62] ), .op(n10775) );
  nand4_1 U11049 ( .ip1(n10778), .ip2(n10777), .ip3(n10776), .ip4(n10775), 
        .op(n10779) );
  nor4_1 U11050 ( .ip1(n10782), .ip2(n10781), .ip3(n10780), .ip4(n10779), .op(
        n11284) );
  nor2_1 U11051 ( .ip1(n11284), .ip2(n10870), .op(n10783) );
  not_ab_or_c_or_d U11052 ( .ip1(n10828), .ip2(n11283), .ip3(n10784), .ip4(
        n10783), .op(n10806) );
  nand2_1 U11053 ( .ip1(n12202), .ip2(\cache_data[7][126] ), .op(n10788) );
  nand2_1 U11054 ( .ip1(n12170), .ip2(\cache_data[11][126] ), .op(n10787) );
  nand2_1 U11055 ( .ip1(n11964), .ip2(\cache_data[0][126] ), .op(n10786) );
  nand2_1 U11056 ( .ip1(n11966), .ip2(\cache_data[10][126] ), .op(n10785) );
  nand4_1 U11057 ( .ip1(n10788), .ip2(n10787), .ip3(n10786), .ip4(n10785), 
        .op(n10804) );
  nand2_1 U11058 ( .ip1(n12241), .ip2(\cache_data[9][126] ), .op(n10792) );
  nand2_1 U11059 ( .ip1(n11965), .ip2(\cache_data[15][126] ), .op(n10791) );
  nand2_1 U11060 ( .ip1(n12234), .ip2(\cache_data[8][126] ), .op(n10790) );
  nand2_1 U11061 ( .ip1(n12164), .ip2(\cache_data[4][126] ), .op(n10789) );
  nand4_1 U11062 ( .ip1(n10792), .ip2(n10791), .ip3(n10790), .ip4(n10789), 
        .op(n10803) );
  nand2_1 U11063 ( .ip1(n11979), .ip2(\cache_data[1][126] ), .op(n10796) );
  nand2_1 U11064 ( .ip1(n11963), .ip2(\cache_data[5][126] ), .op(n10795) );
  nand2_1 U11065 ( .ip1(n12030), .ip2(\cache_data[12][126] ), .op(n10794) );
  nand2_1 U11066 ( .ip1(n11978), .ip2(\cache_data[3][126] ), .op(n10793) );
  nand4_1 U11067 ( .ip1(n10796), .ip2(n10795), .ip3(n10794), .ip4(n10793), 
        .op(n10802) );
  nand2_1 U11068 ( .ip1(n11688), .ip2(\cache_data[14][126] ), .op(n10800) );
  nand2_1 U11069 ( .ip1(n12242), .ip2(\cache_data[13][126] ), .op(n10799) );
  nand2_1 U11070 ( .ip1(n11972), .ip2(\cache_data[6][126] ), .op(n10798) );
  nand2_1 U11071 ( .ip1(n11973), .ip2(\cache_data[2][126] ), .op(n10797) );
  nand4_1 U11072 ( .ip1(n10800), .ip2(n10799), .ip3(n10798), .ip4(n10797), 
        .op(n10801) );
  or4_1 U11073 ( .ip1(n10804), .ip2(n10803), .ip3(n10802), .ip4(n10801), .op(
        n11288) );
  nand2_1 U11074 ( .ip1(n10894), .ip2(n11288), .op(n10805) );
  nand3_1 U11075 ( .ip1(n10807), .ip2(n10806), .ip3(n10805), .op(n7418) );
  nand2_1 U11076 ( .ip1(n12234), .ip2(\cache_data[8][31] ), .op(n10811) );
  nand2_1 U11077 ( .ip1(n12170), .ip2(\cache_data[11][31] ), .op(n10810) );
  nand2_1 U11078 ( .ip1(n11972), .ip2(\cache_data[6][31] ), .op(n10809) );
  nand2_1 U11079 ( .ip1(n12242), .ip2(\cache_data[13][31] ), .op(n10808) );
  nand4_1 U11080 ( .ip1(n10811), .ip2(n10810), .ip3(n10809), .ip4(n10808), 
        .op(n10827) );
  nand2_1 U11081 ( .ip1(n11688), .ip2(\cache_data[14][31] ), .op(n10815) );
  nand2_1 U11082 ( .ip1(n11964), .ip2(\cache_data[0][31] ), .op(n10814) );
  nand2_1 U11083 ( .ip1(n11966), .ip2(\cache_data[10][31] ), .op(n10813) );
  nand2_1 U11084 ( .ip1(n11963), .ip2(\cache_data[5][31] ), .op(n10812) );
  nand4_1 U11085 ( .ip1(n10815), .ip2(n10814), .ip3(n10813), .ip4(n10812), 
        .op(n10826) );
  nand2_1 U11086 ( .ip1(n11943), .ip2(\cache_data[1][31] ), .op(n10819) );
  nand2_1 U11087 ( .ip1(n12030), .ip2(\cache_data[12][31] ), .op(n10818) );
  nand2_1 U11088 ( .ip1(n12164), .ip2(\cache_data[4][31] ), .op(n10817) );
  nand2_1 U11089 ( .ip1(n11973), .ip2(\cache_data[2][31] ), .op(n10816) );
  nand4_1 U11090 ( .ip1(n10819), .ip2(n10818), .ip3(n10817), .ip4(n10816), 
        .op(n10825) );
  nand2_1 U11091 ( .ip1(n12241), .ip2(\cache_data[9][31] ), .op(n10823) );
  nand2_1 U11092 ( .ip1(n12202), .ip2(\cache_data[7][31] ), .op(n10822) );
  nand2_1 U11093 ( .ip1(n11978), .ip2(\cache_data[3][31] ), .op(n10821) );
  nand2_1 U11094 ( .ip1(n11965), .ip2(\cache_data[15][31] ), .op(n10820) );
  nand4_1 U11095 ( .ip1(n10823), .ip2(n10822), .ip3(n10821), .ip4(n10820), 
        .op(n10824) );
  or4_1 U11096 ( .ip1(n10827), .ip2(n10826), .ip3(n10825), .ip4(n10824), .op(
        n11292) );
  nand2_1 U11097 ( .ip1(n10828), .ip2(n11292), .op(n10897) );
  nand2_1 U11098 ( .ip1(n11688), .ip2(\cache_data[14][95] ), .op(n10832) );
  nand2_1 U11099 ( .ip1(n12170), .ip2(\cache_data[11][95] ), .op(n10831) );
  nand2_1 U11100 ( .ip1(n11978), .ip2(\cache_data[3][95] ), .op(n10830) );
  nand2_1 U11101 ( .ip1(n12242), .ip2(\cache_data[13][95] ), .op(n10829) );
  nand4_1 U11102 ( .ip1(n10832), .ip2(n10831), .ip3(n10830), .ip4(n10829), 
        .op(n10848) );
  nand2_1 U11103 ( .ip1(n11943), .ip2(\cache_data[1][95] ), .op(n10836) );
  nand2_1 U11104 ( .ip1(n11965), .ip2(\cache_data[15][95] ), .op(n10835) );
  nand2_1 U11105 ( .ip1(n12234), .ip2(\cache_data[8][95] ), .op(n10834) );
  nand2_1 U11106 ( .ip1(n11972), .ip2(\cache_data[6][95] ), .op(n10833) );
  nand4_1 U11107 ( .ip1(n10836), .ip2(n10835), .ip3(n10834), .ip4(n10833), 
        .op(n10847) );
  nand2_1 U11108 ( .ip1(n11964), .ip2(\cache_data[0][95] ), .op(n10840) );
  nand2_1 U11109 ( .ip1(n12241), .ip2(\cache_data[9][95] ), .op(n10839) );
  nand2_1 U11110 ( .ip1(n11973), .ip2(\cache_data[2][95] ), .op(n10838) );
  nand2_1 U11111 ( .ip1(n12164), .ip2(\cache_data[4][95] ), .op(n10837) );
  nand4_1 U11112 ( .ip1(n10840), .ip2(n10839), .ip3(n10838), .ip4(n10837), 
        .op(n10846) );
  nand2_1 U11113 ( .ip1(n12030), .ip2(\cache_data[12][95] ), .op(n10844) );
  nand2_1 U11114 ( .ip1(n11966), .ip2(\cache_data[10][95] ), .op(n10843) );
  nand2_1 U11115 ( .ip1(n12202), .ip2(\cache_data[7][95] ), .op(n10842) );
  nand2_1 U11116 ( .ip1(n11963), .ip2(\cache_data[5][95] ), .op(n10841) );
  nand4_1 U11117 ( .ip1(n10844), .ip2(n10843), .ip3(n10842), .ip4(n10841), 
        .op(n10845) );
  nor4_1 U11118 ( .ip1(n10848), .ip2(n10847), .ip3(n10846), .ip4(n10845), .op(
        n11295) );
  nor2_1 U11119 ( .ip1(n11295), .ip2(n10849), .op(n10872) );
  nand2_1 U11120 ( .ip1(n11963), .ip2(\cache_data[5][63] ), .op(n10853) );
  nand2_1 U11121 ( .ip1(n11973), .ip2(\cache_data[2][63] ), .op(n10852) );
  nand2_1 U11122 ( .ip1(n11964), .ip2(\cache_data[0][63] ), .op(n10851) );
  nand2_1 U11123 ( .ip1(n11688), .ip2(\cache_data[14][63] ), .op(n10850) );
  nand4_1 U11124 ( .ip1(n10853), .ip2(n10852), .ip3(n10851), .ip4(n10850), 
        .op(n10869) );
  nand2_1 U11125 ( .ip1(n12242), .ip2(\cache_data[13][63] ), .op(n10857) );
  nand2_1 U11126 ( .ip1(n12170), .ip2(\cache_data[11][63] ), .op(n10856) );
  nand2_1 U11127 ( .ip1(n12030), .ip2(\cache_data[12][63] ), .op(n10855) );
  nand2_1 U11128 ( .ip1(n12202), .ip2(\cache_data[7][63] ), .op(n10854) );
  nand4_1 U11129 ( .ip1(n10857), .ip2(n10856), .ip3(n10855), .ip4(n10854), 
        .op(n10868) );
  nand2_1 U11130 ( .ip1(n12234), .ip2(\cache_data[8][63] ), .op(n10861) );
  nand2_1 U11131 ( .ip1(n11966), .ip2(\cache_data[10][63] ), .op(n10860) );
  nand2_1 U11132 ( .ip1(n12241), .ip2(\cache_data[9][63] ), .op(n10859) );
  nand2_1 U11133 ( .ip1(n11979), .ip2(\cache_data[1][63] ), .op(n10858) );
  nand4_1 U11134 ( .ip1(n10861), .ip2(n10860), .ip3(n10859), .ip4(n10858), 
        .op(n10867) );
  nand2_1 U11135 ( .ip1(n12164), .ip2(\cache_data[4][63] ), .op(n10865) );
  nand2_1 U11136 ( .ip1(n11965), .ip2(\cache_data[15][63] ), .op(n10864) );
  nand2_1 U11137 ( .ip1(n11972), .ip2(\cache_data[6][63] ), .op(n10863) );
  nand2_1 U11138 ( .ip1(n11978), .ip2(\cache_data[3][63] ), .op(n10862) );
  nand4_1 U11139 ( .ip1(n10865), .ip2(n10864), .ip3(n10863), .ip4(n10862), 
        .op(n10866) );
  nor4_1 U11140 ( .ip1(n10869), .ip2(n10868), .ip3(n10867), .ip4(n10866), .op(
        n11297) );
  nor2_1 U11141 ( .ip1(n11297), .ip2(n10870), .op(n10871) );
  not_ab_or_c_or_d U11142 ( .ip1(data_wr_mem[31]), .ip2(n10873), .ip3(n10872), 
        .ip4(n10871), .op(n10896) );
  nand2_1 U11143 ( .ip1(n11978), .ip2(\cache_data[3][127] ), .op(n10877) );
  nand2_1 U11144 ( .ip1(n11966), .ip2(\cache_data[10][127] ), .op(n10876) );
  nand2_1 U11145 ( .ip1(n11973), .ip2(\cache_data[2][127] ), .op(n10875) );
  nand2_1 U11146 ( .ip1(n11943), .ip2(\cache_data[1][127] ), .op(n10874) );
  nand4_1 U11147 ( .ip1(n10877), .ip2(n10876), .ip3(n10875), .ip4(n10874), 
        .op(n10893) );
  nand2_1 U11148 ( .ip1(n12241), .ip2(\cache_data[9][127] ), .op(n10881) );
  nand2_1 U11149 ( .ip1(n11688), .ip2(\cache_data[14][127] ), .op(n10880) );
  nand2_1 U11150 ( .ip1(n12202), .ip2(\cache_data[7][127] ), .op(n10879) );
  nand2_1 U11151 ( .ip1(n11972), .ip2(\cache_data[6][127] ), .op(n10878) );
  nand4_1 U11152 ( .ip1(n10881), .ip2(n10880), .ip3(n10879), .ip4(n10878), 
        .op(n10892) );
  nand2_1 U11153 ( .ip1(n12164), .ip2(\cache_data[4][127] ), .op(n10885) );
  nand2_1 U11154 ( .ip1(n11964), .ip2(\cache_data[0][127] ), .op(n10884) );
  nand2_1 U11155 ( .ip1(n12242), .ip2(\cache_data[13][127] ), .op(n10883) );
  nand2_1 U11156 ( .ip1(n11965), .ip2(\cache_data[15][127] ), .op(n10882) );
  nand4_1 U11157 ( .ip1(n10885), .ip2(n10884), .ip3(n10883), .ip4(n10882), 
        .op(n10891) );
  nand2_1 U11158 ( .ip1(n12030), .ip2(\cache_data[12][127] ), .op(n10889) );
  nand2_1 U11159 ( .ip1(n12170), .ip2(\cache_data[11][127] ), .op(n10888) );
  nand2_1 U11160 ( .ip1(n11963), .ip2(\cache_data[5][127] ), .op(n10887) );
  nand2_1 U11161 ( .ip1(n12234), .ip2(\cache_data[8][127] ), .op(n10886) );
  nand4_1 U11162 ( .ip1(n10889), .ip2(n10888), .ip3(n10887), .ip4(n10886), 
        .op(n10890) );
  or4_1 U11163 ( .ip1(n10893), .ip2(n10892), .ip3(n10891), .ip4(n10890), .op(
        n11301) );
  nand2_1 U11164 ( .ip1(n10894), .ip2(n11301), .op(n10895) );
  nand3_1 U11165 ( .ip1(n10897), .ip2(n10896), .ip3(n10895), .op(n7417) );
  nand2_1 U11166 ( .ip1(n10898), .ip2(n12325), .op(n10977) );
  nand2_1 U11167 ( .ip1(n12252), .ip2(n10977), .op(n11658) );
  and2_1 U11168 ( .ip1(n11658), .ip2(mem_data_cnt[2]), .op(n10899) );
  xor2_1 U11169 ( .ip1(mem_data_cnt[3]), .ip2(n10899), .op(n7416) );
  mux2_1 U11170 ( .ip1(mem_data_cnt[2]), .ip2(n11433), .s(n11658), .op(n7415)
         );
  inv_1 U11171 ( .ip(n12323), .op(n11307) );
  nand2_1 U11172 ( .ip1(n11307), .ip2(n10900), .op(n12257) );
  nand2_1 U11173 ( .ip1(wr_mem), .ip2(n12257), .op(n10901) );
  nand2_1 U11174 ( .ip1(n12252), .ip2(n10901), .op(n7414) );
  nand2_1 U11175 ( .ip1(rd_mem), .ip2(n12257), .op(n10902) );
  nand2_1 U11176 ( .ip1(n10977), .ip2(n10902), .op(n7413) );
  nand2_1 U11177 ( .ip1(cache_valid[7]), .ip2(n10933), .op(n10920) );
  nand2_1 U11178 ( .ip1(n10949), .ip2(cache_valid[13]), .op(n10905) );
  nand2_1 U11179 ( .ip1(n10924), .ip2(cache_valid[6]), .op(n10904) );
  nand2_1 U11180 ( .ip1(n10922), .ip2(cache_valid[10]), .op(n10903) );
  nand3_1 U11181 ( .ip1(n10905), .ip2(n10904), .ip3(n10903), .op(n10915) );
  and2_1 U11182 ( .ip1(n10947), .ip2(cache_valid[5]), .op(n10907) );
  and2_1 U11183 ( .ip1(n10923), .ip2(cache_valid[9]), .op(n10906) );
  not_ab_or_c_or_d U11184 ( .ip1(cache_valid[2]), .ip2(n10925), .ip3(n10907), 
        .ip4(n10906), .op(n10913) );
  and2_1 U11185 ( .ip1(n10930), .ip2(cache_valid[1]), .op(n10909) );
  and2_1 U11186 ( .ip1(n10941), .ip2(cache_valid[11]), .op(n10908) );
  not_ab_or_c_or_d U11187 ( .ip1(cache_valid[14]), .ip2(n10938), .ip3(n10909), 
        .ip4(n10908), .op(n10912) );
  nand2_1 U11188 ( .ip1(n10931), .ip2(cache_valid[3]), .op(n10911) );
  nand2_1 U11189 ( .ip1(n10939), .ip2(cache_valid[12]), .op(n10910) );
  nand4_1 U11190 ( .ip1(n10913), .ip2(n10912), .ip3(n10911), .ip4(n10910), 
        .op(n10914) );
  not_ab_or_c_or_d U11191 ( .ip1(n10948), .ip2(cache_valid[4]), .ip3(n10915), 
        .ip4(n10914), .op(n10919) );
  and2_1 U11192 ( .ip1(n10932), .ip2(cache_valid[8]), .op(n10917) );
  and2_1 U11193 ( .ip1(n10940), .ip2(cache_valid[15]), .op(n10916) );
  not_ab_or_c_or_d U11194 ( .ip1(cache_valid[0]), .ip2(n10946), .ip3(n10917), 
        .ip4(n10916), .op(n10918) );
  nand3_1 U11195 ( .ip1(n10920), .ip2(n10919), .ip3(n10918), .op(n10921) );
  mux2_1 U11196 ( .ip1(valid), .ip2(n10921), .s(n11358), .op(n7411) );
  nand2_1 U11197 ( .ip1(n10922), .ip2(cache_dirty[10]), .op(n10929) );
  nand2_1 U11198 ( .ip1(n10923), .ip2(cache_dirty[9]), .op(n10928) );
  nand2_1 U11199 ( .ip1(n10924), .ip2(cache_dirty[6]), .op(n10927) );
  nand2_1 U11200 ( .ip1(n10925), .ip2(cache_dirty[2]), .op(n10926) );
  nand4_1 U11201 ( .ip1(n10929), .ip2(n10928), .ip3(n10927), .ip4(n10926), 
        .op(n10957) );
  nand2_1 U11202 ( .ip1(n10930), .ip2(cache_dirty[1]), .op(n10937) );
  nand2_1 U11203 ( .ip1(n10931), .ip2(cache_dirty[3]), .op(n10936) );
  nand2_1 U11204 ( .ip1(n10932), .ip2(cache_dirty[8]), .op(n10935) );
  nand2_1 U11205 ( .ip1(n10933), .ip2(cache_dirty[7]), .op(n10934) );
  nand4_1 U11206 ( .ip1(n10937), .ip2(n10936), .ip3(n10935), .ip4(n10934), 
        .op(n10956) );
  nand2_1 U11207 ( .ip1(n10938), .ip2(cache_dirty[14]), .op(n10945) );
  nand2_1 U11208 ( .ip1(n10939), .ip2(cache_dirty[12]), .op(n10944) );
  nand2_1 U11209 ( .ip1(n10940), .ip2(cache_dirty[15]), .op(n10943) );
  nand2_1 U11210 ( .ip1(n10941), .ip2(cache_dirty[11]), .op(n10942) );
  nand4_1 U11211 ( .ip1(n10945), .ip2(n10944), .ip3(n10943), .ip4(n10942), 
        .op(n10955) );
  nand2_1 U11212 ( .ip1(n10946), .ip2(cache_dirty[0]), .op(n10953) );
  nand2_1 U11213 ( .ip1(n10947), .ip2(cache_dirty[5]), .op(n10952) );
  nand2_1 U11214 ( .ip1(n10948), .ip2(cache_dirty[4]), .op(n10951) );
  nand2_1 U11215 ( .ip1(n10949), .ip2(cache_dirty[13]), .op(n10950) );
  nand4_1 U11216 ( .ip1(n10953), .ip2(n10952), .ip3(n10951), .ip4(n10950), 
        .op(n10954) );
  or4_1 U11217 ( .ip1(n10957), .ip2(n10956), .ip3(n10955), .ip4(n10954), .op(
        n10958) );
  mux2_1 U11218 ( .ip1(dirty), .ip2(n10958), .s(n11358), .op(n7410) );
  mux2_1 U11219 ( .ip1(N3615), .ip2(addr_req[0]), .s(n11358), .op(n7409) );
  and2_1 U11220 ( .ip1(n11361), .ip2(N3616), .op(n7408) );
  mux2_1 U11221 ( .ip1(N3612), .ip2(addr_req[1]), .s(n11358), .op(n7407) );
  and2_1 U11222 ( .ip1(n11361), .ip2(N3613), .op(n7406) );
  mux2_1 U11223 ( .ip1(N3609), .ip2(addr_req[2]), .s(n11358), .op(n7405) );
  and2_1 U11224 ( .ip1(n11361), .ip2(N3610), .op(n7404) );
  mux2_1 U11225 ( .ip1(N3606), .ip2(addr_req[3]), .s(n11358), .op(n7403) );
  and2_1 U11226 ( .ip1(n11361), .ip2(N3607), .op(n7402) );
  mux2_1 U11227 ( .ip1(N3603), .ip2(addr_req[4]), .s(n11358), .op(n7401) );
  and2_1 U11228 ( .ip1(n11361), .ip2(N3604), .op(n7400) );
  mux2_1 U11229 ( .ip1(N3600), .ip2(addr_req[5]), .s(n11358), .op(n7399) );
  and2_1 U11230 ( .ip1(n11361), .ip2(N3601), .op(n7398) );
  mux2_1 U11231 ( .ip1(N3597), .ip2(addr_req[6]), .s(n7728), .op(n7397) );
  and2_1 U11232 ( .ip1(n11361), .ip2(N3598), .op(n7396) );
  mux2_1 U11233 ( .ip1(N3594), .ip2(addr_req[7]), .s(n7728), .op(n7395) );
  and2_1 U11234 ( .ip1(n11361), .ip2(N3595), .op(n7394) );
  inv_1 U11235 ( .ip(n10977), .op(n12254) );
  nand2_1 U11236 ( .ip1(n12233), .ip2(n12254), .op(n11308) );
  inv_1 U11237 ( .ip(cache_valid[0]), .op(n10959) );
  nand2_1 U11238 ( .ip1(n11308), .ip2(n10959), .op(n7393) );
  nand2_1 U11239 ( .ip1(n11979), .ip2(n12254), .op(n11311) );
  inv_1 U11240 ( .ip(cache_valid[1]), .op(n10960) );
  nand2_1 U11241 ( .ip1(n11311), .ip2(n10960), .op(n7392) );
  nand2_1 U11242 ( .ip1(n11973), .ip2(n12254), .op(n11314) );
  inv_1 U11243 ( .ip(cache_valid[2]), .op(n10961) );
  nand2_1 U11244 ( .ip1(n11314), .ip2(n10961), .op(n7391) );
  nand2_1 U11245 ( .ip1(n11978), .ip2(n12254), .op(n11318) );
  inv_1 U11246 ( .ip(cache_valid[3]), .op(n10962) );
  nand2_1 U11247 ( .ip1(n11318), .ip2(n10962), .op(n7390) );
  nand2_1 U11248 ( .ip1(n12164), .ip2(n12254), .op(n11321) );
  inv_1 U11249 ( .ip(cache_valid[4]), .op(n10963) );
  nand2_1 U11250 ( .ip1(n11321), .ip2(n10963), .op(n7389) );
  nand2_1 U11251 ( .ip1(n10964), .ip2(n12254), .op(n11324) );
  inv_1 U11252 ( .ip(cache_valid[5]), .op(n10965) );
  nand2_1 U11253 ( .ip1(n11324), .ip2(n10965), .op(n7388) );
  nand2_1 U11254 ( .ip1(n11972), .ip2(n12254), .op(n11327) );
  inv_1 U11255 ( .ip(cache_valid[6]), .op(n10966) );
  nand2_1 U11256 ( .ip1(n11327), .ip2(n10966), .op(n7387) );
  nand2_1 U11257 ( .ip1(n12202), .ip2(n12254), .op(n11330) );
  inv_1 U11258 ( .ip(cache_valid[7]), .op(n10967) );
  nand2_1 U11259 ( .ip1(n11330), .ip2(n10967), .op(n7386) );
  nand2_1 U11260 ( .ip1(n12234), .ip2(n12254), .op(n11333) );
  inv_1 U11261 ( .ip(cache_valid[8]), .op(n10968) );
  nand2_1 U11262 ( .ip1(n11333), .ip2(n10968), .op(n7385) );
  nand2_1 U11263 ( .ip1(n12241), .ip2(n12254), .op(n11336) );
  inv_1 U11264 ( .ip(cache_valid[9]), .op(n10969) );
  nand2_1 U11265 ( .ip1(n11336), .ip2(n10969), .op(n7384) );
  nand2_1 U11266 ( .ip1(n12196), .ip2(n12254), .op(n11339) );
  inv_1 U11267 ( .ip(cache_valid[10]), .op(n10970) );
  nand2_1 U11268 ( .ip1(n11339), .ip2(n10970), .op(n7383) );
  nand2_1 U11269 ( .ip1(n12170), .ip2(n12254), .op(n11342) );
  inv_1 U11270 ( .ip(cache_valid[11]), .op(n10971) );
  nand2_1 U11271 ( .ip1(n11342), .ip2(n10971), .op(n7382) );
  nand2_1 U11272 ( .ip1(n12030), .ip2(n12254), .op(n11345) );
  inv_1 U11273 ( .ip(cache_valid[12]), .op(n10972) );
  nand2_1 U11274 ( .ip1(n11345), .ip2(n10972), .op(n7381) );
  nand2_1 U11275 ( .ip1(n12242), .ip2(n12254), .op(n11348) );
  inv_1 U11276 ( .ip(cache_valid[13]), .op(n10973) );
  nand2_1 U11277 ( .ip1(n11348), .ip2(n10973), .op(n7380) );
  nand2_1 U11278 ( .ip1(n11688), .ip2(n12254), .op(n11351) );
  inv_1 U11279 ( .ip(cache_valid[14]), .op(n10974) );
  nand2_1 U11280 ( .ip1(n11351), .ip2(n10974), .op(n7379) );
  nand2_1 U11281 ( .ip1(n10975), .ip2(n12254), .op(n11354) );
  inv_1 U11282 ( .ip(cache_valid[15]), .op(n10976) );
  nand2_1 U11283 ( .ip1(n11354), .ip2(n10976), .op(n7378) );
  mux2_1 U11284 ( .ip1(N3591), .ip2(addr_req[8]), .s(n7728), .op(n7377) );
  and2_1 U11285 ( .ip1(n11361), .ip2(N3592), .op(n7376) );
  nor3_1 U11286 ( .ip1(n12324), .ip2(n8923), .ip3(n10977), .op(n10994) );
  buf_1 U11287 ( .ip(n10994), .op(n10978) );
  mux2_1 U11288 ( .ip1(\cache_tag[0][0] ), .ip2(addr_resp[8]), .s(n10978), 
        .op(n7375) );
  nor3_1 U11289 ( .ip1(n12324), .ip2(n11459), .ip3(n10977), .op(n10995) );
  buf_1 U11290 ( .ip(n10995), .op(n10979) );
  mux2_1 U11291 ( .ip1(\cache_tag[1][0] ), .ip2(addr_resp[8]), .s(n10979), 
        .op(n7374) );
  nor3_1 U11292 ( .ip1(n12324), .ip2(n8928), .ip3(n10977), .op(n10996) );
  buf_1 U11293 ( .ip(n10996), .op(n10980) );
  mux2_1 U11294 ( .ip1(\cache_tag[2][0] ), .ip2(addr_resp[8]), .s(n10980), 
        .op(n7373) );
  nor3_1 U11295 ( .ip1(n12324), .ip2(n11476), .ip3(n10977), .op(n10997) );
  buf_1 U11296 ( .ip(n10997), .op(n10981) );
  mux2_1 U11297 ( .ip1(\cache_tag[3][0] ), .ip2(addr_resp[8]), .s(n10981), 
        .op(n7372) );
  nor3_1 U11298 ( .ip1(n12324), .ip2(n8136), .ip3(n10977), .op(n10998) );
  buf_1 U11299 ( .ip(n10998), .op(n10982) );
  mux2_1 U11300 ( .ip1(\cache_tag[4][0] ), .ip2(addr_resp[8]), .s(n10982), 
        .op(n7371) );
  nor3_1 U11301 ( .ip1(n12324), .ip2(n11493), .ip3(n10977), .op(n10999) );
  buf_1 U11302 ( .ip(n10999), .op(n10983) );
  mux2_1 U11303 ( .ip1(\cache_tag[5][0] ), .ip2(addr_resp[8]), .s(n10983), 
        .op(n7370) );
  nor3_1 U11304 ( .ip1(n12324), .ip2(n11502), .ip3(n10977), .op(n11000) );
  buf_1 U11305 ( .ip(n11000), .op(n10984) );
  mux2_1 U11306 ( .ip1(\cache_tag[6][0] ), .ip2(addr_resp[8]), .s(n10984), 
        .op(n7369) );
  nor3_1 U11307 ( .ip1(n12324), .ip2(n8153), .ip3(n10977), .op(n11001) );
  buf_1 U11308 ( .ip(n11001), .op(n10985) );
  mux2_1 U11309 ( .ip1(\cache_tag[7][0] ), .ip2(addr_resp[8]), .s(n10985), 
        .op(n7368) );
  nor3_1 U11310 ( .ip1(n12324), .ip2(n8137), .ip3(n10977), .op(n11002) );
  buf_1 U11311 ( .ip(n11002), .op(n10986) );
  mux2_1 U11312 ( .ip1(\cache_tag[8][0] ), .ip2(addr_resp[8]), .s(n10986), 
        .op(n7367) );
  nor3_1 U11313 ( .ip1(n12324), .ip2(n8144), .ip3(n10977), .op(n11003) );
  buf_1 U11314 ( .ip(n11003), .op(n10987) );
  mux2_1 U11315 ( .ip1(\cache_tag[9][0] ), .ip2(addr_resp[8]), .s(n10987), 
        .op(n7366) );
  nor3_1 U11316 ( .ip1(n12324), .ip2(n8146), .ip3(n10977), .op(n11004) );
  buf_1 U11317 ( .ip(n11004), .op(n10988) );
  mux2_1 U11318 ( .ip1(\cache_tag[10][0] ), .ip2(addr_resp[8]), .s(n10988), 
        .op(n7365) );
  nor3_1 U11319 ( .ip1(n12324), .ip2(n8151), .ip3(n10977), .op(n11005) );
  buf_1 U11320 ( .ip(n11005), .op(n10989) );
  mux2_1 U11321 ( .ip1(\cache_tag[11][0] ), .ip2(addr_resp[8]), .s(n10989), 
        .op(n7364) );
  inv_1 U11322 ( .ip(n12030), .op(n11551) );
  nor3_1 U11323 ( .ip1(n12324), .ip2(n11551), .ip3(n10977), .op(n11006) );
  buf_1 U11324 ( .ip(n11006), .op(n10990) );
  mux2_1 U11325 ( .ip1(\cache_tag[12][0] ), .ip2(addr_resp[8]), .s(n10990), 
        .op(n7363) );
  nor3_1 U11326 ( .ip1(rst), .ip2(n8145), .ip3(n10977), .op(n11007) );
  buf_1 U11327 ( .ip(n11007), .op(n10991) );
  mux2_1 U11328 ( .ip1(\cache_tag[13][0] ), .ip2(addr_resp[8]), .s(n10991), 
        .op(n7362) );
  nor3_1 U11329 ( .ip1(rst), .ip2(n11600), .ip3(n10977), .op(n11008) );
  buf_1 U11330 ( .ip(n11008), .op(n10992) );
  mux2_1 U11331 ( .ip1(\cache_tag[14][0] ), .ip2(addr_resp[8]), .s(n10992), 
        .op(n7361) );
  nor3_1 U11332 ( .ip1(n12324), .ip2(n11612), .ip3(n10977), .op(n11009) );
  buf_1 U11333 ( .ip(n11009), .op(n10993) );
  mux2_1 U11334 ( .ip1(\cache_tag[15][0] ), .ip2(addr_resp[8]), .s(n10993), 
        .op(n7360) );
  mux2_1 U11335 ( .ip1(N3588), .ip2(addr_req[9]), .s(n7728), .op(n7359) );
  and2_1 U11336 ( .ip1(n11361), .ip2(N3589), .op(n7358) );
  mux2_1 U11337 ( .ip1(\cache_tag[0][1] ), .ip2(addr_resp[9]), .s(n10978), 
        .op(n7357) );
  mux2_1 U11338 ( .ip1(\cache_tag[1][1] ), .ip2(addr_resp[9]), .s(n10979), 
        .op(n7356) );
  mux2_1 U11339 ( .ip1(\cache_tag[2][1] ), .ip2(addr_resp[9]), .s(n10980), 
        .op(n7355) );
  mux2_1 U11340 ( .ip1(\cache_tag[3][1] ), .ip2(addr_resp[9]), .s(n10981), 
        .op(n7354) );
  mux2_1 U11341 ( .ip1(\cache_tag[4][1] ), .ip2(addr_resp[9]), .s(n10982), 
        .op(n7353) );
  mux2_1 U11342 ( .ip1(\cache_tag[5][1] ), .ip2(addr_resp[9]), .s(n10983), 
        .op(n7352) );
  mux2_1 U11343 ( .ip1(\cache_tag[6][1] ), .ip2(addr_resp[9]), .s(n10984), 
        .op(n7351) );
  mux2_1 U11344 ( .ip1(\cache_tag[7][1] ), .ip2(addr_resp[9]), .s(n10985), 
        .op(n7350) );
  mux2_1 U11345 ( .ip1(\cache_tag[8][1] ), .ip2(addr_resp[9]), .s(n10986), 
        .op(n7349) );
  mux2_1 U11346 ( .ip1(\cache_tag[9][1] ), .ip2(addr_resp[9]), .s(n10987), 
        .op(n7348) );
  mux2_1 U11347 ( .ip1(\cache_tag[10][1] ), .ip2(addr_resp[9]), .s(n10988), 
        .op(n7347) );
  mux2_1 U11348 ( .ip1(\cache_tag[11][1] ), .ip2(addr_resp[9]), .s(n10989), 
        .op(n7346) );
  mux2_1 U11349 ( .ip1(\cache_tag[12][1] ), .ip2(addr_resp[9]), .s(n10990), 
        .op(n7345) );
  mux2_1 U11350 ( .ip1(\cache_tag[13][1] ), .ip2(addr_resp[9]), .s(n10991), 
        .op(n7344) );
  mux2_1 U11351 ( .ip1(\cache_tag[14][1] ), .ip2(addr_resp[9]), .s(n10992), 
        .op(n7343) );
  mux2_1 U11352 ( .ip1(\cache_tag[15][1] ), .ip2(addr_resp[9]), .s(n10993), 
        .op(n7342) );
  mux2_1 U11353 ( .ip1(N3585), .ip2(addr_req[10]), .s(n7728), .op(n7341) );
  and2_1 U11354 ( .ip1(n11361), .ip2(N3586), .op(n7340) );
  mux2_1 U11355 ( .ip1(\cache_tag[0][2] ), .ip2(addr_resp[10]), .s(n10978), 
        .op(n7339) );
  mux2_1 U11356 ( .ip1(\cache_tag[1][2] ), .ip2(addr_resp[10]), .s(n10979), 
        .op(n7338) );
  mux2_1 U11357 ( .ip1(\cache_tag[2][2] ), .ip2(addr_resp[10]), .s(n10980), 
        .op(n7337) );
  mux2_1 U11358 ( .ip1(\cache_tag[3][2] ), .ip2(addr_resp[10]), .s(n10981), 
        .op(n7336) );
  mux2_1 U11359 ( .ip1(\cache_tag[4][2] ), .ip2(addr_resp[10]), .s(n10982), 
        .op(n7335) );
  mux2_1 U11360 ( .ip1(\cache_tag[5][2] ), .ip2(addr_resp[10]), .s(n10983), 
        .op(n7334) );
  mux2_1 U11361 ( .ip1(\cache_tag[6][2] ), .ip2(addr_resp[10]), .s(n10984), 
        .op(n7333) );
  mux2_1 U11362 ( .ip1(\cache_tag[7][2] ), .ip2(addr_resp[10]), .s(n10985), 
        .op(n7332) );
  mux2_1 U11363 ( .ip1(\cache_tag[8][2] ), .ip2(addr_resp[10]), .s(n10986), 
        .op(n7331) );
  mux2_1 U11364 ( .ip1(\cache_tag[9][2] ), .ip2(addr_resp[10]), .s(n10987), 
        .op(n7330) );
  mux2_1 U11365 ( .ip1(\cache_tag[10][2] ), .ip2(addr_resp[10]), .s(n10988), 
        .op(n7329) );
  mux2_1 U11366 ( .ip1(\cache_tag[11][2] ), .ip2(addr_resp[10]), .s(n10989), 
        .op(n7328) );
  mux2_1 U11367 ( .ip1(\cache_tag[12][2] ), .ip2(addr_resp[10]), .s(n10990), 
        .op(n7327) );
  mux2_1 U11368 ( .ip1(\cache_tag[13][2] ), .ip2(addr_resp[10]), .s(n10991), 
        .op(n7326) );
  mux2_1 U11369 ( .ip1(\cache_tag[14][2] ), .ip2(addr_resp[10]), .s(n10992), 
        .op(n7325) );
  mux2_1 U11370 ( .ip1(\cache_tag[15][2] ), .ip2(addr_resp[10]), .s(n10993), 
        .op(n7324) );
  mux2_1 U11371 ( .ip1(N3582), .ip2(addr_req[11]), .s(n7728), .op(n7323) );
  and2_1 U11372 ( .ip1(n11361), .ip2(N3583), .op(n7322) );
  mux2_1 U11373 ( .ip1(\cache_tag[0][3] ), .ip2(addr_resp[11]), .s(n10978), 
        .op(n7321) );
  mux2_1 U11374 ( .ip1(\cache_tag[1][3] ), .ip2(addr_resp[11]), .s(n10979), 
        .op(n7320) );
  mux2_1 U11375 ( .ip1(\cache_tag[2][3] ), .ip2(addr_resp[11]), .s(n10980), 
        .op(n7319) );
  mux2_1 U11376 ( .ip1(\cache_tag[3][3] ), .ip2(addr_resp[11]), .s(n10981), 
        .op(n7318) );
  mux2_1 U11377 ( .ip1(\cache_tag[4][3] ), .ip2(addr_resp[11]), .s(n10982), 
        .op(n7317) );
  mux2_1 U11378 ( .ip1(\cache_tag[5][3] ), .ip2(addr_resp[11]), .s(n10983), 
        .op(n7316) );
  mux2_1 U11379 ( .ip1(\cache_tag[6][3] ), .ip2(addr_resp[11]), .s(n10984), 
        .op(n7315) );
  mux2_1 U11380 ( .ip1(\cache_tag[7][3] ), .ip2(addr_resp[11]), .s(n10985), 
        .op(n7314) );
  mux2_1 U11381 ( .ip1(\cache_tag[8][3] ), .ip2(addr_resp[11]), .s(n10986), 
        .op(n7313) );
  mux2_1 U11382 ( .ip1(\cache_tag[9][3] ), .ip2(addr_resp[11]), .s(n10987), 
        .op(n7312) );
  mux2_1 U11383 ( .ip1(\cache_tag[10][3] ), .ip2(addr_resp[11]), .s(n10988), 
        .op(n7311) );
  mux2_1 U11384 ( .ip1(\cache_tag[11][3] ), .ip2(addr_resp[11]), .s(n10989), 
        .op(n7310) );
  mux2_1 U11385 ( .ip1(\cache_tag[12][3] ), .ip2(addr_resp[11]), .s(n10990), 
        .op(n7309) );
  mux2_1 U11386 ( .ip1(\cache_tag[13][3] ), .ip2(addr_resp[11]), .s(n10991), 
        .op(n7308) );
  mux2_1 U11387 ( .ip1(\cache_tag[14][3] ), .ip2(addr_resp[11]), .s(n10992), 
        .op(n7307) );
  mux2_1 U11388 ( .ip1(\cache_tag[15][3] ), .ip2(addr_resp[11]), .s(n10993), 
        .op(n7306) );
  mux2_1 U11389 ( .ip1(N3579), .ip2(addr_req[12]), .s(n7728), .op(n7305) );
  and2_1 U11390 ( .ip1(n11361), .ip2(N3580), .op(n7304) );
  mux2_1 U11391 ( .ip1(\cache_tag[0][4] ), .ip2(addr_resp[12]), .s(n10978), 
        .op(n7303) );
  mux2_1 U11392 ( .ip1(\cache_tag[1][4] ), .ip2(addr_resp[12]), .s(n10979), 
        .op(n7302) );
  mux2_1 U11393 ( .ip1(\cache_tag[2][4] ), .ip2(addr_resp[12]), .s(n10980), 
        .op(n7301) );
  mux2_1 U11394 ( .ip1(\cache_tag[3][4] ), .ip2(addr_resp[12]), .s(n10981), 
        .op(n7300) );
  mux2_1 U11395 ( .ip1(\cache_tag[4][4] ), .ip2(addr_resp[12]), .s(n10982), 
        .op(n7299) );
  mux2_1 U11396 ( .ip1(\cache_tag[5][4] ), .ip2(addr_resp[12]), .s(n10983), 
        .op(n7298) );
  mux2_1 U11397 ( .ip1(\cache_tag[6][4] ), .ip2(addr_resp[12]), .s(n10984), 
        .op(n7297) );
  mux2_1 U11398 ( .ip1(\cache_tag[7][4] ), .ip2(addr_resp[12]), .s(n10985), 
        .op(n7296) );
  mux2_1 U11399 ( .ip1(\cache_tag[8][4] ), .ip2(addr_resp[12]), .s(n10986), 
        .op(n7295) );
  mux2_1 U11400 ( .ip1(\cache_tag[9][4] ), .ip2(addr_resp[12]), .s(n10987), 
        .op(n7294) );
  mux2_1 U11401 ( .ip1(\cache_tag[10][4] ), .ip2(addr_resp[12]), .s(n10988), 
        .op(n7293) );
  mux2_1 U11402 ( .ip1(\cache_tag[11][4] ), .ip2(addr_resp[12]), .s(n10989), 
        .op(n7292) );
  mux2_1 U11403 ( .ip1(\cache_tag[12][4] ), .ip2(addr_resp[12]), .s(n10990), 
        .op(n7291) );
  mux2_1 U11404 ( .ip1(\cache_tag[13][4] ), .ip2(addr_resp[12]), .s(n10991), 
        .op(n7290) );
  mux2_1 U11405 ( .ip1(\cache_tag[14][4] ), .ip2(addr_resp[12]), .s(n10992), 
        .op(n7289) );
  mux2_1 U11406 ( .ip1(\cache_tag[15][4] ), .ip2(addr_resp[12]), .s(n10993), 
        .op(n7288) );
  mux2_1 U11407 ( .ip1(N3576), .ip2(addr_req[13]), .s(n7728), .op(n7287) );
  and2_1 U11408 ( .ip1(n11361), .ip2(N3577), .op(n7286) );
  mux2_1 U11409 ( .ip1(\cache_tag[0][5] ), .ip2(addr_resp[13]), .s(n10978), 
        .op(n7285) );
  mux2_1 U11410 ( .ip1(\cache_tag[1][5] ), .ip2(addr_resp[13]), .s(n10979), 
        .op(n7284) );
  mux2_1 U11411 ( .ip1(\cache_tag[2][5] ), .ip2(addr_resp[13]), .s(n10980), 
        .op(n7283) );
  mux2_1 U11412 ( .ip1(\cache_tag[3][5] ), .ip2(addr_resp[13]), .s(n10981), 
        .op(n7282) );
  mux2_1 U11413 ( .ip1(\cache_tag[4][5] ), .ip2(addr_resp[13]), .s(n10982), 
        .op(n7281) );
  mux2_1 U11414 ( .ip1(\cache_tag[5][5] ), .ip2(addr_resp[13]), .s(n10983), 
        .op(n7280) );
  mux2_1 U11415 ( .ip1(\cache_tag[6][5] ), .ip2(addr_resp[13]), .s(n10984), 
        .op(n7279) );
  mux2_1 U11416 ( .ip1(\cache_tag[7][5] ), .ip2(addr_resp[13]), .s(n10985), 
        .op(n7278) );
  mux2_1 U11417 ( .ip1(\cache_tag[8][5] ), .ip2(addr_resp[13]), .s(n10986), 
        .op(n7277) );
  mux2_1 U11418 ( .ip1(\cache_tag[9][5] ), .ip2(addr_resp[13]), .s(n10987), 
        .op(n7276) );
  mux2_1 U11419 ( .ip1(\cache_tag[10][5] ), .ip2(addr_resp[13]), .s(n10988), 
        .op(n7275) );
  mux2_1 U11420 ( .ip1(\cache_tag[11][5] ), .ip2(addr_resp[13]), .s(n10989), 
        .op(n7274) );
  mux2_1 U11421 ( .ip1(\cache_tag[12][5] ), .ip2(addr_resp[13]), .s(n10990), 
        .op(n7273) );
  mux2_1 U11422 ( .ip1(\cache_tag[13][5] ), .ip2(addr_resp[13]), .s(n10991), 
        .op(n7272) );
  mux2_1 U11423 ( .ip1(\cache_tag[14][5] ), .ip2(addr_resp[13]), .s(n10992), 
        .op(n7271) );
  mux2_1 U11424 ( .ip1(\cache_tag[15][5] ), .ip2(addr_resp[13]), .s(n10993), 
        .op(n7270) );
  mux2_1 U11425 ( .ip1(N3573), .ip2(addr_req[14]), .s(n7728), .op(n7269) );
  and2_1 U11426 ( .ip1(n11361), .ip2(N3574), .op(n7268) );
  mux2_1 U11427 ( .ip1(\cache_tag[0][6] ), .ip2(addr_resp[14]), .s(n10978), 
        .op(n7267) );
  mux2_1 U11428 ( .ip1(\cache_tag[1][6] ), .ip2(addr_resp[14]), .s(n10979), 
        .op(n7266) );
  mux2_1 U11429 ( .ip1(\cache_tag[2][6] ), .ip2(addr_resp[14]), .s(n10980), 
        .op(n7265) );
  mux2_1 U11430 ( .ip1(\cache_tag[3][6] ), .ip2(addr_resp[14]), .s(n10981), 
        .op(n7264) );
  mux2_1 U11431 ( .ip1(\cache_tag[4][6] ), .ip2(addr_resp[14]), .s(n10982), 
        .op(n7263) );
  mux2_1 U11432 ( .ip1(\cache_tag[5][6] ), .ip2(addr_resp[14]), .s(n10983), 
        .op(n7262) );
  mux2_1 U11433 ( .ip1(\cache_tag[6][6] ), .ip2(addr_resp[14]), .s(n10984), 
        .op(n7261) );
  mux2_1 U11434 ( .ip1(\cache_tag[7][6] ), .ip2(addr_resp[14]), .s(n10985), 
        .op(n7260) );
  mux2_1 U11435 ( .ip1(\cache_tag[8][6] ), .ip2(addr_resp[14]), .s(n10986), 
        .op(n7259) );
  mux2_1 U11436 ( .ip1(\cache_tag[9][6] ), .ip2(addr_resp[14]), .s(n10987), 
        .op(n7258) );
  mux2_1 U11437 ( .ip1(\cache_tag[10][6] ), .ip2(addr_resp[14]), .s(n10988), 
        .op(n7257) );
  mux2_1 U11438 ( .ip1(\cache_tag[11][6] ), .ip2(addr_resp[14]), .s(n10989), 
        .op(n7256) );
  mux2_1 U11439 ( .ip1(\cache_tag[12][6] ), .ip2(addr_resp[14]), .s(n10990), 
        .op(n7255) );
  mux2_1 U11440 ( .ip1(\cache_tag[13][6] ), .ip2(addr_resp[14]), .s(n10991), 
        .op(n7254) );
  mux2_1 U11441 ( .ip1(\cache_tag[14][6] ), .ip2(addr_resp[14]), .s(n10992), 
        .op(n7253) );
  mux2_1 U11442 ( .ip1(\cache_tag[15][6] ), .ip2(addr_resp[14]), .s(n10993), 
        .op(n7252) );
  mux2_1 U11443 ( .ip1(N3570), .ip2(addr_req[15]), .s(n7728), .op(n7251) );
  and2_1 U11444 ( .ip1(n11361), .ip2(N3571), .op(n7250) );
  mux2_1 U11445 ( .ip1(\cache_tag[0][7] ), .ip2(addr_resp[15]), .s(n10978), 
        .op(n7249) );
  mux2_1 U11446 ( .ip1(\cache_tag[1][7] ), .ip2(addr_resp[15]), .s(n10979), 
        .op(n7248) );
  mux2_1 U11447 ( .ip1(\cache_tag[2][7] ), .ip2(addr_resp[15]), .s(n10980), 
        .op(n7247) );
  mux2_1 U11448 ( .ip1(\cache_tag[3][7] ), .ip2(addr_resp[15]), .s(n10981), 
        .op(n7246) );
  mux2_1 U11449 ( .ip1(\cache_tag[4][7] ), .ip2(addr_resp[15]), .s(n10982), 
        .op(n7245) );
  mux2_1 U11450 ( .ip1(\cache_tag[5][7] ), .ip2(addr_resp[15]), .s(n10983), 
        .op(n7244) );
  mux2_1 U11451 ( .ip1(\cache_tag[6][7] ), .ip2(addr_resp[15]), .s(n10984), 
        .op(n7243) );
  mux2_1 U11452 ( .ip1(\cache_tag[7][7] ), .ip2(addr_resp[15]), .s(n10985), 
        .op(n7242) );
  mux2_1 U11453 ( .ip1(\cache_tag[8][7] ), .ip2(addr_resp[15]), .s(n10986), 
        .op(n7241) );
  mux2_1 U11454 ( .ip1(\cache_tag[9][7] ), .ip2(addr_resp[15]), .s(n10987), 
        .op(n7240) );
  mux2_1 U11455 ( .ip1(\cache_tag[10][7] ), .ip2(addr_resp[15]), .s(n10988), 
        .op(n7239) );
  mux2_1 U11456 ( .ip1(\cache_tag[11][7] ), .ip2(addr_resp[15]), .s(n10989), 
        .op(n7238) );
  mux2_1 U11457 ( .ip1(\cache_tag[12][7] ), .ip2(addr_resp[15]), .s(n10990), 
        .op(n7237) );
  mux2_1 U11458 ( .ip1(\cache_tag[13][7] ), .ip2(addr_resp[15]), .s(n10991), 
        .op(n7236) );
  mux2_1 U11459 ( .ip1(\cache_tag[14][7] ), .ip2(addr_resp[15]), .s(n10992), 
        .op(n7235) );
  mux2_1 U11460 ( .ip1(\cache_tag[15][7] ), .ip2(addr_resp[15]), .s(n10993), 
        .op(n7234) );
  mux2_1 U11461 ( .ip1(N3567), .ip2(addr_req[16]), .s(n11358), .op(n7233) );
  and2_1 U11462 ( .ip1(n11361), .ip2(N3568), .op(n7232) );
  mux2_1 U11463 ( .ip1(\cache_tag[0][8] ), .ip2(addr_resp[16]), .s(n10978), 
        .op(n7231) );
  mux2_1 U11464 ( .ip1(\cache_tag[1][8] ), .ip2(addr_resp[16]), .s(n10979), 
        .op(n7230) );
  mux2_1 U11465 ( .ip1(\cache_tag[2][8] ), .ip2(addr_resp[16]), .s(n10980), 
        .op(n7229) );
  mux2_1 U11466 ( .ip1(\cache_tag[3][8] ), .ip2(addr_resp[16]), .s(n10981), 
        .op(n7228) );
  mux2_1 U11467 ( .ip1(\cache_tag[4][8] ), .ip2(addr_resp[16]), .s(n10982), 
        .op(n7227) );
  mux2_1 U11468 ( .ip1(\cache_tag[5][8] ), .ip2(addr_resp[16]), .s(n10983), 
        .op(n7226) );
  mux2_1 U11469 ( .ip1(\cache_tag[6][8] ), .ip2(addr_resp[16]), .s(n10984), 
        .op(n7225) );
  mux2_1 U11470 ( .ip1(\cache_tag[7][8] ), .ip2(addr_resp[16]), .s(n10985), 
        .op(n7224) );
  mux2_1 U11471 ( .ip1(\cache_tag[8][8] ), .ip2(addr_resp[16]), .s(n10986), 
        .op(n7223) );
  mux2_1 U11472 ( .ip1(\cache_tag[9][8] ), .ip2(addr_resp[16]), .s(n10987), 
        .op(n7222) );
  mux2_1 U11473 ( .ip1(\cache_tag[10][8] ), .ip2(addr_resp[16]), .s(n10988), 
        .op(n7221) );
  mux2_1 U11474 ( .ip1(\cache_tag[11][8] ), .ip2(addr_resp[16]), .s(n10989), 
        .op(n7220) );
  mux2_1 U11475 ( .ip1(\cache_tag[12][8] ), .ip2(addr_resp[16]), .s(n10990), 
        .op(n7219) );
  mux2_1 U11476 ( .ip1(\cache_tag[13][8] ), .ip2(addr_resp[16]), .s(n10991), 
        .op(n7218) );
  mux2_1 U11477 ( .ip1(\cache_tag[14][8] ), .ip2(addr_resp[16]), .s(n10992), 
        .op(n7217) );
  mux2_1 U11478 ( .ip1(\cache_tag[15][8] ), .ip2(addr_resp[16]), .s(n10993), 
        .op(n7216) );
  mux2_1 U11479 ( .ip1(N3564), .ip2(addr_req[17]), .s(n11358), .op(n7215) );
  and2_1 U11480 ( .ip1(n11361), .ip2(N3565), .op(n7214) );
  mux2_1 U11481 ( .ip1(\cache_tag[0][9] ), .ip2(addr_resp[17]), .s(n10978), 
        .op(n7213) );
  mux2_1 U11482 ( .ip1(\cache_tag[1][9] ), .ip2(addr_resp[17]), .s(n10979), 
        .op(n7212) );
  mux2_1 U11483 ( .ip1(\cache_tag[2][9] ), .ip2(addr_resp[17]), .s(n10980), 
        .op(n7211) );
  mux2_1 U11484 ( .ip1(\cache_tag[3][9] ), .ip2(addr_resp[17]), .s(n10981), 
        .op(n7210) );
  mux2_1 U11485 ( .ip1(\cache_tag[4][9] ), .ip2(addr_resp[17]), .s(n10982), 
        .op(n7209) );
  mux2_1 U11486 ( .ip1(\cache_tag[5][9] ), .ip2(addr_resp[17]), .s(n10983), 
        .op(n7208) );
  mux2_1 U11487 ( .ip1(\cache_tag[6][9] ), .ip2(addr_resp[17]), .s(n10984), 
        .op(n7207) );
  mux2_1 U11488 ( .ip1(\cache_tag[7][9] ), .ip2(addr_resp[17]), .s(n10985), 
        .op(n7206) );
  mux2_1 U11489 ( .ip1(\cache_tag[8][9] ), .ip2(addr_resp[17]), .s(n10986), 
        .op(n7205) );
  mux2_1 U11490 ( .ip1(\cache_tag[9][9] ), .ip2(addr_resp[17]), .s(n10987), 
        .op(n7204) );
  mux2_1 U11491 ( .ip1(\cache_tag[10][9] ), .ip2(addr_resp[17]), .s(n10988), 
        .op(n7203) );
  mux2_1 U11492 ( .ip1(\cache_tag[11][9] ), .ip2(addr_resp[17]), .s(n10989), 
        .op(n7202) );
  mux2_1 U11493 ( .ip1(\cache_tag[12][9] ), .ip2(addr_resp[17]), .s(n10990), 
        .op(n7201) );
  mux2_1 U11494 ( .ip1(\cache_tag[13][9] ), .ip2(addr_resp[17]), .s(n10991), 
        .op(n7200) );
  mux2_1 U11495 ( .ip1(\cache_tag[14][9] ), .ip2(addr_resp[17]), .s(n10992), 
        .op(n7199) );
  mux2_1 U11496 ( .ip1(\cache_tag[15][9] ), .ip2(addr_resp[17]), .s(n10993), 
        .op(n7198) );
  mux2_1 U11497 ( .ip1(N3561), .ip2(addr_req[18]), .s(n11358), .op(n7197) );
  and2_1 U11498 ( .ip1(n11361), .ip2(N3562), .op(n7196) );
  mux2_1 U11499 ( .ip1(\cache_tag[0][10] ), .ip2(addr_resp[18]), .s(n10978), 
        .op(n7195) );
  mux2_1 U11500 ( .ip1(\cache_tag[1][10] ), .ip2(addr_resp[18]), .s(n10979), 
        .op(n7194) );
  mux2_1 U11501 ( .ip1(\cache_tag[2][10] ), .ip2(addr_resp[18]), .s(n10980), 
        .op(n7193) );
  mux2_1 U11502 ( .ip1(\cache_tag[3][10] ), .ip2(addr_resp[18]), .s(n10981), 
        .op(n7192) );
  mux2_1 U11503 ( .ip1(\cache_tag[4][10] ), .ip2(addr_resp[18]), .s(n10982), 
        .op(n7191) );
  mux2_1 U11504 ( .ip1(\cache_tag[5][10] ), .ip2(addr_resp[18]), .s(n10983), 
        .op(n7190) );
  mux2_1 U11505 ( .ip1(\cache_tag[6][10] ), .ip2(addr_resp[18]), .s(n10984), 
        .op(n7189) );
  mux2_1 U11506 ( .ip1(\cache_tag[7][10] ), .ip2(addr_resp[18]), .s(n10985), 
        .op(n7188) );
  mux2_1 U11507 ( .ip1(\cache_tag[8][10] ), .ip2(addr_resp[18]), .s(n10986), 
        .op(n7187) );
  mux2_1 U11508 ( .ip1(\cache_tag[9][10] ), .ip2(addr_resp[18]), .s(n10987), 
        .op(n7186) );
  mux2_1 U11509 ( .ip1(\cache_tag[10][10] ), .ip2(addr_resp[18]), .s(n10988), 
        .op(n7185) );
  mux2_1 U11510 ( .ip1(\cache_tag[11][10] ), .ip2(addr_resp[18]), .s(n10989), 
        .op(n7184) );
  mux2_1 U11511 ( .ip1(\cache_tag[12][10] ), .ip2(addr_resp[18]), .s(n10990), 
        .op(n7183) );
  mux2_1 U11512 ( .ip1(\cache_tag[13][10] ), .ip2(addr_resp[18]), .s(n10991), 
        .op(n7182) );
  mux2_1 U11513 ( .ip1(\cache_tag[14][10] ), .ip2(addr_resp[18]), .s(n10992), 
        .op(n7181) );
  mux2_1 U11514 ( .ip1(\cache_tag[15][10] ), .ip2(addr_resp[18]), .s(n10993), 
        .op(n7180) );
  mux2_1 U11515 ( .ip1(N3558), .ip2(addr_req[19]), .s(n7728), .op(n7179) );
  and2_1 U11516 ( .ip1(n11361), .ip2(N3559), .op(n7178) );
  mux2_1 U11517 ( .ip1(\cache_tag[0][11] ), .ip2(addr_resp[19]), .s(n10978), 
        .op(n7177) );
  mux2_1 U11518 ( .ip1(\cache_tag[1][11] ), .ip2(addr_resp[19]), .s(n10979), 
        .op(n7176) );
  mux2_1 U11519 ( .ip1(\cache_tag[2][11] ), .ip2(addr_resp[19]), .s(n10980), 
        .op(n7175) );
  mux2_1 U11520 ( .ip1(\cache_tag[3][11] ), .ip2(addr_resp[19]), .s(n10981), 
        .op(n7174) );
  mux2_1 U11521 ( .ip1(\cache_tag[4][11] ), .ip2(addr_resp[19]), .s(n10982), 
        .op(n7173) );
  mux2_1 U11522 ( .ip1(\cache_tag[5][11] ), .ip2(addr_resp[19]), .s(n10983), 
        .op(n7172) );
  mux2_1 U11523 ( .ip1(\cache_tag[6][11] ), .ip2(addr_resp[19]), .s(n10984), 
        .op(n7171) );
  mux2_1 U11524 ( .ip1(\cache_tag[7][11] ), .ip2(addr_resp[19]), .s(n10985), 
        .op(n7170) );
  mux2_1 U11525 ( .ip1(\cache_tag[8][11] ), .ip2(addr_resp[19]), .s(n10986), 
        .op(n7169) );
  mux2_1 U11526 ( .ip1(\cache_tag[9][11] ), .ip2(addr_resp[19]), .s(n10987), 
        .op(n7168) );
  mux2_1 U11527 ( .ip1(\cache_tag[10][11] ), .ip2(addr_resp[19]), .s(n10988), 
        .op(n7167) );
  mux2_1 U11528 ( .ip1(\cache_tag[11][11] ), .ip2(addr_resp[19]), .s(n10989), 
        .op(n7166) );
  mux2_1 U11529 ( .ip1(\cache_tag[12][11] ), .ip2(addr_resp[19]), .s(n10990), 
        .op(n7165) );
  mux2_1 U11530 ( .ip1(\cache_tag[13][11] ), .ip2(addr_resp[19]), .s(n10991), 
        .op(n7164) );
  mux2_1 U11531 ( .ip1(\cache_tag[14][11] ), .ip2(addr_resp[19]), .s(n10992), 
        .op(n7163) );
  mux2_1 U11532 ( .ip1(\cache_tag[15][11] ), .ip2(addr_resp[19]), .s(n10993), 
        .op(n7162) );
  mux2_1 U11533 ( .ip1(N3555), .ip2(addr_req[20]), .s(n7728), .op(n7161) );
  and2_1 U11534 ( .ip1(n11361), .ip2(N3556), .op(n7160) );
  mux2_1 U11535 ( .ip1(\cache_tag[0][12] ), .ip2(addr_resp[20]), .s(n10978), 
        .op(n7159) );
  mux2_1 U11536 ( .ip1(\cache_tag[1][12] ), .ip2(addr_resp[20]), .s(n10979), 
        .op(n7158) );
  mux2_1 U11537 ( .ip1(\cache_tag[2][12] ), .ip2(addr_resp[20]), .s(n10980), 
        .op(n7157) );
  mux2_1 U11538 ( .ip1(\cache_tag[3][12] ), .ip2(addr_resp[20]), .s(n10981), 
        .op(n7156) );
  mux2_1 U11539 ( .ip1(\cache_tag[4][12] ), .ip2(addr_resp[20]), .s(n10982), 
        .op(n7155) );
  mux2_1 U11540 ( .ip1(\cache_tag[5][12] ), .ip2(addr_resp[20]), .s(n10983), 
        .op(n7154) );
  mux2_1 U11541 ( .ip1(\cache_tag[6][12] ), .ip2(addr_resp[20]), .s(n10984), 
        .op(n7153) );
  mux2_1 U11542 ( .ip1(\cache_tag[7][12] ), .ip2(addr_resp[20]), .s(n10985), 
        .op(n7152) );
  mux2_1 U11543 ( .ip1(\cache_tag[8][12] ), .ip2(addr_resp[20]), .s(n10986), 
        .op(n7151) );
  mux2_1 U11544 ( .ip1(\cache_tag[9][12] ), .ip2(addr_resp[20]), .s(n10987), 
        .op(n7150) );
  mux2_1 U11545 ( .ip1(\cache_tag[10][12] ), .ip2(addr_resp[20]), .s(n10988), 
        .op(n7149) );
  mux2_1 U11546 ( .ip1(\cache_tag[11][12] ), .ip2(addr_resp[20]), .s(n10989), 
        .op(n7148) );
  mux2_1 U11547 ( .ip1(\cache_tag[12][12] ), .ip2(addr_resp[20]), .s(n10990), 
        .op(n7147) );
  mux2_1 U11548 ( .ip1(\cache_tag[13][12] ), .ip2(addr_resp[20]), .s(n10991), 
        .op(n7146) );
  mux2_1 U11549 ( .ip1(\cache_tag[14][12] ), .ip2(addr_resp[20]), .s(n10992), 
        .op(n7145) );
  mux2_1 U11550 ( .ip1(\cache_tag[15][12] ), .ip2(addr_resp[20]), .s(n10993), 
        .op(n7144) );
  mux2_1 U11551 ( .ip1(N3552), .ip2(addr_req[21]), .s(n7728), .op(n7143) );
  and2_1 U11552 ( .ip1(n11361), .ip2(N3553), .op(n7142) );
  mux2_1 U11553 ( .ip1(\cache_tag[0][13] ), .ip2(addr_resp[21]), .s(n10978), 
        .op(n7141) );
  mux2_1 U11554 ( .ip1(\cache_tag[1][13] ), .ip2(addr_resp[21]), .s(n10979), 
        .op(n7140) );
  mux2_1 U11555 ( .ip1(\cache_tag[2][13] ), .ip2(addr_resp[21]), .s(n10980), 
        .op(n7139) );
  mux2_1 U11556 ( .ip1(\cache_tag[3][13] ), .ip2(addr_resp[21]), .s(n10981), 
        .op(n7138) );
  mux2_1 U11557 ( .ip1(\cache_tag[4][13] ), .ip2(addr_resp[21]), .s(n10982), 
        .op(n7137) );
  mux2_1 U11558 ( .ip1(\cache_tag[5][13] ), .ip2(addr_resp[21]), .s(n10983), 
        .op(n7136) );
  mux2_1 U11559 ( .ip1(\cache_tag[6][13] ), .ip2(addr_resp[21]), .s(n10984), 
        .op(n7135) );
  mux2_1 U11560 ( .ip1(\cache_tag[7][13] ), .ip2(addr_resp[21]), .s(n10985), 
        .op(n7134) );
  mux2_1 U11561 ( .ip1(\cache_tag[8][13] ), .ip2(addr_resp[21]), .s(n10986), 
        .op(n7133) );
  mux2_1 U11562 ( .ip1(\cache_tag[9][13] ), .ip2(addr_resp[21]), .s(n10987), 
        .op(n7132) );
  mux2_1 U11563 ( .ip1(\cache_tag[10][13] ), .ip2(addr_resp[21]), .s(n10988), 
        .op(n7131) );
  mux2_1 U11564 ( .ip1(\cache_tag[11][13] ), .ip2(addr_resp[21]), .s(n10989), 
        .op(n7130) );
  mux2_1 U11565 ( .ip1(\cache_tag[12][13] ), .ip2(addr_resp[21]), .s(n10990), 
        .op(n7129) );
  mux2_1 U11566 ( .ip1(\cache_tag[13][13] ), .ip2(addr_resp[21]), .s(n10991), 
        .op(n7128) );
  mux2_1 U11567 ( .ip1(\cache_tag[14][13] ), .ip2(addr_resp[21]), .s(n10992), 
        .op(n7127) );
  mux2_1 U11568 ( .ip1(\cache_tag[15][13] ), .ip2(addr_resp[21]), .s(n10993), 
        .op(n7126) );
  mux2_1 U11569 ( .ip1(N3549), .ip2(addr_req[22]), .s(n7728), .op(n7125) );
  and2_1 U11570 ( .ip1(n11361), .ip2(N3550), .op(n7124) );
  mux2_1 U11571 ( .ip1(\cache_tag[0][14] ), .ip2(addr_resp[22]), .s(n10978), 
        .op(n7123) );
  mux2_1 U11572 ( .ip1(\cache_tag[1][14] ), .ip2(addr_resp[22]), .s(n10979), 
        .op(n7122) );
  mux2_1 U11573 ( .ip1(\cache_tag[2][14] ), .ip2(addr_resp[22]), .s(n10980), 
        .op(n7121) );
  mux2_1 U11574 ( .ip1(\cache_tag[3][14] ), .ip2(addr_resp[22]), .s(n10981), 
        .op(n7120) );
  mux2_1 U11575 ( .ip1(\cache_tag[4][14] ), .ip2(addr_resp[22]), .s(n10982), 
        .op(n7119) );
  mux2_1 U11576 ( .ip1(\cache_tag[5][14] ), .ip2(addr_resp[22]), .s(n10983), 
        .op(n7118) );
  mux2_1 U11577 ( .ip1(\cache_tag[6][14] ), .ip2(addr_resp[22]), .s(n10984), 
        .op(n7117) );
  mux2_1 U11578 ( .ip1(\cache_tag[7][14] ), .ip2(addr_resp[22]), .s(n10985), 
        .op(n7116) );
  mux2_1 U11579 ( .ip1(\cache_tag[8][14] ), .ip2(addr_resp[22]), .s(n10986), 
        .op(n7115) );
  mux2_1 U11580 ( .ip1(\cache_tag[9][14] ), .ip2(addr_resp[22]), .s(n10987), 
        .op(n7114) );
  mux2_1 U11581 ( .ip1(\cache_tag[10][14] ), .ip2(addr_resp[22]), .s(n10988), 
        .op(n7113) );
  mux2_1 U11582 ( .ip1(\cache_tag[11][14] ), .ip2(addr_resp[22]), .s(n10989), 
        .op(n7112) );
  mux2_1 U11583 ( .ip1(\cache_tag[12][14] ), .ip2(addr_resp[22]), .s(n10990), 
        .op(n7111) );
  mux2_1 U11584 ( .ip1(\cache_tag[13][14] ), .ip2(addr_resp[22]), .s(n10991), 
        .op(n7110) );
  mux2_1 U11585 ( .ip1(\cache_tag[14][14] ), .ip2(addr_resp[22]), .s(n10992), 
        .op(n7109) );
  mux2_1 U11586 ( .ip1(\cache_tag[15][14] ), .ip2(addr_resp[22]), .s(n10993), 
        .op(n7108) );
  mux2_1 U11587 ( .ip1(N3546), .ip2(addr_req[23]), .s(n7728), .op(n7107) );
  and2_1 U11588 ( .ip1(n11361), .ip2(N3547), .op(n7106) );
  mux2_1 U11589 ( .ip1(\cache_tag[0][15] ), .ip2(addr_resp[23]), .s(n10978), 
        .op(n7105) );
  mux2_1 U11590 ( .ip1(\cache_tag[1][15] ), .ip2(addr_resp[23]), .s(n10979), 
        .op(n7104) );
  mux2_1 U11591 ( .ip1(\cache_tag[2][15] ), .ip2(addr_resp[23]), .s(n10980), 
        .op(n7103) );
  mux2_1 U11592 ( .ip1(\cache_tag[3][15] ), .ip2(addr_resp[23]), .s(n10981), 
        .op(n7102) );
  mux2_1 U11593 ( .ip1(\cache_tag[4][15] ), .ip2(addr_resp[23]), .s(n10982), 
        .op(n7101) );
  mux2_1 U11594 ( .ip1(\cache_tag[5][15] ), .ip2(addr_resp[23]), .s(n10983), 
        .op(n7100) );
  mux2_1 U11595 ( .ip1(\cache_tag[6][15] ), .ip2(addr_resp[23]), .s(n10984), 
        .op(n7099) );
  mux2_1 U11596 ( .ip1(\cache_tag[7][15] ), .ip2(addr_resp[23]), .s(n10985), 
        .op(n7098) );
  mux2_1 U11597 ( .ip1(\cache_tag[8][15] ), .ip2(addr_resp[23]), .s(n10986), 
        .op(n7097) );
  mux2_1 U11598 ( .ip1(\cache_tag[9][15] ), .ip2(addr_resp[23]), .s(n10987), 
        .op(n7096) );
  mux2_1 U11599 ( .ip1(\cache_tag[10][15] ), .ip2(addr_resp[23]), .s(n10988), 
        .op(n7095) );
  mux2_1 U11600 ( .ip1(\cache_tag[11][15] ), .ip2(addr_resp[23]), .s(n10989), 
        .op(n7094) );
  mux2_1 U11601 ( .ip1(\cache_tag[12][15] ), .ip2(addr_resp[23]), .s(n10990), 
        .op(n7093) );
  mux2_1 U11602 ( .ip1(\cache_tag[13][15] ), .ip2(addr_resp[23]), .s(n10991), 
        .op(n7092) );
  mux2_1 U11603 ( .ip1(\cache_tag[14][15] ), .ip2(addr_resp[23]), .s(n10992), 
        .op(n7091) );
  mux2_1 U11604 ( .ip1(\cache_tag[15][15] ), .ip2(addr_resp[23]), .s(n10993), 
        .op(n7090) );
  mux2_1 U11605 ( .ip1(N3543), .ip2(addr_req[24]), .s(n11358), .op(n7089) );
  and2_1 U11606 ( .ip1(n11361), .ip2(N3544), .op(n7088) );
  mux2_1 U11607 ( .ip1(\cache_tag[0][16] ), .ip2(addr_resp[24]), .s(n10994), 
        .op(n7087) );
  mux2_1 U11608 ( .ip1(\cache_tag[1][16] ), .ip2(addr_resp[24]), .s(n10995), 
        .op(n7086) );
  mux2_1 U11609 ( .ip1(\cache_tag[2][16] ), .ip2(addr_resp[24]), .s(n10996), 
        .op(n7085) );
  mux2_1 U11610 ( .ip1(\cache_tag[3][16] ), .ip2(addr_resp[24]), .s(n10997), 
        .op(n7084) );
  mux2_1 U11611 ( .ip1(\cache_tag[4][16] ), .ip2(addr_resp[24]), .s(n10998), 
        .op(n7083) );
  mux2_1 U11612 ( .ip1(\cache_tag[5][16] ), .ip2(addr_resp[24]), .s(n10999), 
        .op(n7082) );
  mux2_1 U11613 ( .ip1(\cache_tag[6][16] ), .ip2(addr_resp[24]), .s(n11000), 
        .op(n7081) );
  mux2_1 U11614 ( .ip1(\cache_tag[7][16] ), .ip2(addr_resp[24]), .s(n11001), 
        .op(n7080) );
  mux2_1 U11615 ( .ip1(\cache_tag[8][16] ), .ip2(addr_resp[24]), .s(n11002), 
        .op(n7079) );
  mux2_1 U11616 ( .ip1(\cache_tag[9][16] ), .ip2(addr_resp[24]), .s(n11003), 
        .op(n7078) );
  mux2_1 U11617 ( .ip1(\cache_tag[10][16] ), .ip2(addr_resp[24]), .s(n11004), 
        .op(n7077) );
  mux2_1 U11618 ( .ip1(\cache_tag[11][16] ), .ip2(addr_resp[24]), .s(n11005), 
        .op(n7076) );
  mux2_1 U11619 ( .ip1(\cache_tag[12][16] ), .ip2(addr_resp[24]), .s(n11006), 
        .op(n7075) );
  mux2_1 U11620 ( .ip1(\cache_tag[13][16] ), .ip2(addr_resp[24]), .s(n11007), 
        .op(n7074) );
  mux2_1 U11621 ( .ip1(\cache_tag[14][16] ), .ip2(addr_resp[24]), .s(n11008), 
        .op(n7073) );
  mux2_1 U11622 ( .ip1(\cache_tag[15][16] ), .ip2(addr_resp[24]), .s(n11009), 
        .op(n7072) );
  mux2_1 U11623 ( .ip1(N3540), .ip2(addr_req[25]), .s(n7728), .op(n7071) );
  and2_1 U11624 ( .ip1(n11361), .ip2(N3541), .op(n7070) );
  mux2_1 U11625 ( .ip1(\cache_tag[0][17] ), .ip2(addr_resp[25]), .s(n10994), 
        .op(n7069) );
  mux2_1 U11626 ( .ip1(\cache_tag[1][17] ), .ip2(addr_resp[25]), .s(n10995), 
        .op(n7068) );
  mux2_1 U11627 ( .ip1(\cache_tag[2][17] ), .ip2(addr_resp[25]), .s(n10996), 
        .op(n7067) );
  mux2_1 U11628 ( .ip1(\cache_tag[3][17] ), .ip2(addr_resp[25]), .s(n10997), 
        .op(n7066) );
  mux2_1 U11629 ( .ip1(\cache_tag[4][17] ), .ip2(addr_resp[25]), .s(n10998), 
        .op(n7065) );
  mux2_1 U11630 ( .ip1(\cache_tag[5][17] ), .ip2(addr_resp[25]), .s(n10999), 
        .op(n7064) );
  mux2_1 U11631 ( .ip1(\cache_tag[6][17] ), .ip2(addr_resp[25]), .s(n11000), 
        .op(n7063) );
  mux2_1 U11632 ( .ip1(\cache_tag[7][17] ), .ip2(addr_resp[25]), .s(n11001), 
        .op(n7062) );
  mux2_1 U11633 ( .ip1(\cache_tag[8][17] ), .ip2(addr_resp[25]), .s(n11002), 
        .op(n7061) );
  mux2_1 U11634 ( .ip1(\cache_tag[9][17] ), .ip2(addr_resp[25]), .s(n11003), 
        .op(n7060) );
  mux2_1 U11635 ( .ip1(\cache_tag[10][17] ), .ip2(addr_resp[25]), .s(n11004), 
        .op(n7059) );
  mux2_1 U11636 ( .ip1(\cache_tag[11][17] ), .ip2(addr_resp[25]), .s(n11005), 
        .op(n7058) );
  mux2_1 U11637 ( .ip1(\cache_tag[12][17] ), .ip2(addr_resp[25]), .s(n11006), 
        .op(n7057) );
  mux2_1 U11638 ( .ip1(\cache_tag[13][17] ), .ip2(addr_resp[25]), .s(n11007), 
        .op(n7056) );
  mux2_1 U11639 ( .ip1(\cache_tag[14][17] ), .ip2(addr_resp[25]), .s(n11008), 
        .op(n7055) );
  mux2_1 U11640 ( .ip1(\cache_tag[15][17] ), .ip2(addr_resp[25]), .s(n11009), 
        .op(n7054) );
  mux2_1 U11641 ( .ip1(N3537), .ip2(addr_req[26]), .s(n7728), .op(n7053) );
  and2_1 U11642 ( .ip1(n11361), .ip2(N3538), .op(n7052) );
  mux2_1 U11643 ( .ip1(\cache_tag[0][18] ), .ip2(addr_resp[26]), .s(n10994), 
        .op(n7051) );
  mux2_1 U11644 ( .ip1(\cache_tag[1][18] ), .ip2(addr_resp[26]), .s(n10995), 
        .op(n7050) );
  mux2_1 U11645 ( .ip1(\cache_tag[2][18] ), .ip2(addr_resp[26]), .s(n10996), 
        .op(n7049) );
  mux2_1 U11646 ( .ip1(\cache_tag[3][18] ), .ip2(addr_resp[26]), .s(n10997), 
        .op(n7048) );
  mux2_1 U11647 ( .ip1(\cache_tag[4][18] ), .ip2(addr_resp[26]), .s(n10998), 
        .op(n7047) );
  mux2_1 U11648 ( .ip1(\cache_tag[5][18] ), .ip2(addr_resp[26]), .s(n10999), 
        .op(n7046) );
  mux2_1 U11649 ( .ip1(\cache_tag[6][18] ), .ip2(addr_resp[26]), .s(n11000), 
        .op(n7045) );
  mux2_1 U11650 ( .ip1(\cache_tag[7][18] ), .ip2(addr_resp[26]), .s(n11001), 
        .op(n7044) );
  mux2_1 U11651 ( .ip1(\cache_tag[8][18] ), .ip2(addr_resp[26]), .s(n11002), 
        .op(n7043) );
  mux2_1 U11652 ( .ip1(\cache_tag[9][18] ), .ip2(addr_resp[26]), .s(n11003), 
        .op(n7042) );
  mux2_1 U11653 ( .ip1(\cache_tag[10][18] ), .ip2(addr_resp[26]), .s(n11004), 
        .op(n7041) );
  mux2_1 U11654 ( .ip1(\cache_tag[11][18] ), .ip2(addr_resp[26]), .s(n11005), 
        .op(n7040) );
  mux2_1 U11655 ( .ip1(\cache_tag[12][18] ), .ip2(addr_resp[26]), .s(n11006), 
        .op(n7039) );
  mux2_1 U11656 ( .ip1(\cache_tag[13][18] ), .ip2(addr_resp[26]), .s(n11007), 
        .op(n7038) );
  mux2_1 U11657 ( .ip1(\cache_tag[14][18] ), .ip2(addr_resp[26]), .s(n11008), 
        .op(n7037) );
  mux2_1 U11658 ( .ip1(\cache_tag[15][18] ), .ip2(addr_resp[26]), .s(n11009), 
        .op(n7036) );
  mux2_1 U11659 ( .ip1(N3534), .ip2(addr_req[27]), .s(n7728), .op(n7035) );
  and2_1 U11660 ( .ip1(n11361), .ip2(N3535), .op(n7034) );
  mux2_1 U11661 ( .ip1(\cache_tag[0][19] ), .ip2(addr_resp[27]), .s(n10994), 
        .op(n7033) );
  mux2_1 U11662 ( .ip1(\cache_tag[1][19] ), .ip2(addr_resp[27]), .s(n10995), 
        .op(n7032) );
  mux2_1 U11663 ( .ip1(\cache_tag[2][19] ), .ip2(addr_resp[27]), .s(n10996), 
        .op(n7031) );
  mux2_1 U11664 ( .ip1(\cache_tag[3][19] ), .ip2(addr_resp[27]), .s(n10997), 
        .op(n7030) );
  mux2_1 U11665 ( .ip1(\cache_tag[4][19] ), .ip2(addr_resp[27]), .s(n10998), 
        .op(n7029) );
  mux2_1 U11666 ( .ip1(\cache_tag[5][19] ), .ip2(addr_resp[27]), .s(n10999), 
        .op(n7028) );
  mux2_1 U11667 ( .ip1(\cache_tag[6][19] ), .ip2(addr_resp[27]), .s(n11000), 
        .op(n7027) );
  mux2_1 U11668 ( .ip1(\cache_tag[7][19] ), .ip2(addr_resp[27]), .s(n11001), 
        .op(n7026) );
  mux2_1 U11669 ( .ip1(\cache_tag[8][19] ), .ip2(addr_resp[27]), .s(n11002), 
        .op(n7025) );
  mux2_1 U11670 ( .ip1(\cache_tag[9][19] ), .ip2(addr_resp[27]), .s(n11003), 
        .op(n7024) );
  mux2_1 U11671 ( .ip1(\cache_tag[10][19] ), .ip2(addr_resp[27]), .s(n11004), 
        .op(n7023) );
  mux2_1 U11672 ( .ip1(\cache_tag[11][19] ), .ip2(addr_resp[27]), .s(n11005), 
        .op(n7022) );
  mux2_1 U11673 ( .ip1(\cache_tag[12][19] ), .ip2(addr_resp[27]), .s(n11006), 
        .op(n7021) );
  mux2_1 U11674 ( .ip1(\cache_tag[13][19] ), .ip2(addr_resp[27]), .s(n11007), 
        .op(n7020) );
  mux2_1 U11675 ( .ip1(\cache_tag[14][19] ), .ip2(addr_resp[27]), .s(n11008), 
        .op(n7019) );
  mux2_1 U11676 ( .ip1(\cache_tag[15][19] ), .ip2(addr_resp[27]), .s(n11009), 
        .op(n7018) );
  mux2_1 U11677 ( .ip1(N3531), .ip2(addr_req[28]), .s(n11358), .op(n7017) );
  and2_1 U11678 ( .ip1(n11361), .ip2(N3532), .op(n7016) );
  mux2_1 U11679 ( .ip1(\cache_tag[0][20] ), .ip2(addr_resp[28]), .s(n10994), 
        .op(n7015) );
  mux2_1 U11680 ( .ip1(\cache_tag[1][20] ), .ip2(addr_resp[28]), .s(n10995), 
        .op(n7014) );
  mux2_1 U11681 ( .ip1(\cache_tag[2][20] ), .ip2(addr_resp[28]), .s(n10996), 
        .op(n7013) );
  mux2_1 U11682 ( .ip1(\cache_tag[3][20] ), .ip2(addr_resp[28]), .s(n10997), 
        .op(n7012) );
  mux2_1 U11683 ( .ip1(\cache_tag[4][20] ), .ip2(addr_resp[28]), .s(n10998), 
        .op(n7011) );
  mux2_1 U11684 ( .ip1(\cache_tag[5][20] ), .ip2(addr_resp[28]), .s(n10999), 
        .op(n7010) );
  mux2_1 U11685 ( .ip1(\cache_tag[6][20] ), .ip2(addr_resp[28]), .s(n11000), 
        .op(n7009) );
  mux2_1 U11686 ( .ip1(\cache_tag[7][20] ), .ip2(addr_resp[28]), .s(n11001), 
        .op(n7008) );
  mux2_1 U11687 ( .ip1(\cache_tag[8][20] ), .ip2(addr_resp[28]), .s(n11002), 
        .op(n7007) );
  mux2_1 U11688 ( .ip1(\cache_tag[9][20] ), .ip2(addr_resp[28]), .s(n11003), 
        .op(n7006) );
  mux2_1 U11689 ( .ip1(\cache_tag[10][20] ), .ip2(addr_resp[28]), .s(n11004), 
        .op(n7005) );
  mux2_1 U11690 ( .ip1(\cache_tag[11][20] ), .ip2(addr_resp[28]), .s(n11005), 
        .op(n7004) );
  mux2_1 U11691 ( .ip1(\cache_tag[12][20] ), .ip2(addr_resp[28]), .s(n11006), 
        .op(n7003) );
  mux2_1 U11692 ( .ip1(\cache_tag[13][20] ), .ip2(addr_resp[28]), .s(n11007), 
        .op(n7002) );
  mux2_1 U11693 ( .ip1(\cache_tag[14][20] ), .ip2(addr_resp[28]), .s(n11008), 
        .op(n7001) );
  mux2_1 U11694 ( .ip1(\cache_tag[15][20] ), .ip2(addr_resp[28]), .s(n11009), 
        .op(n7000) );
  mux2_1 U11695 ( .ip1(N3528), .ip2(addr_req[29]), .s(n7728), .op(n6999) );
  and2_1 U11696 ( .ip1(n11361), .ip2(N3529), .op(n6998) );
  mux2_1 U11697 ( .ip1(\cache_tag[0][21] ), .ip2(addr_resp[29]), .s(n10994), 
        .op(n6997) );
  mux2_1 U11698 ( .ip1(\cache_tag[1][21] ), .ip2(addr_resp[29]), .s(n10995), 
        .op(n6996) );
  mux2_1 U11699 ( .ip1(\cache_tag[2][21] ), .ip2(addr_resp[29]), .s(n10996), 
        .op(n6995) );
  mux2_1 U11700 ( .ip1(\cache_tag[3][21] ), .ip2(addr_resp[29]), .s(n10997), 
        .op(n6994) );
  mux2_1 U11701 ( .ip1(\cache_tag[4][21] ), .ip2(addr_resp[29]), .s(n10998), 
        .op(n6993) );
  mux2_1 U11702 ( .ip1(\cache_tag[5][21] ), .ip2(addr_resp[29]), .s(n10999), 
        .op(n6992) );
  mux2_1 U11703 ( .ip1(\cache_tag[6][21] ), .ip2(addr_resp[29]), .s(n11000), 
        .op(n6991) );
  mux2_1 U11704 ( .ip1(\cache_tag[7][21] ), .ip2(addr_resp[29]), .s(n11001), 
        .op(n6990) );
  mux2_1 U11705 ( .ip1(\cache_tag[8][21] ), .ip2(addr_resp[29]), .s(n11002), 
        .op(n6989) );
  mux2_1 U11706 ( .ip1(\cache_tag[9][21] ), .ip2(addr_resp[29]), .s(n11003), 
        .op(n6988) );
  mux2_1 U11707 ( .ip1(\cache_tag[10][21] ), .ip2(addr_resp[29]), .s(n11004), 
        .op(n6987) );
  mux2_1 U11708 ( .ip1(\cache_tag[11][21] ), .ip2(addr_resp[29]), .s(n11005), 
        .op(n6986) );
  mux2_1 U11709 ( .ip1(\cache_tag[12][21] ), .ip2(addr_resp[29]), .s(n11006), 
        .op(n6985) );
  mux2_1 U11710 ( .ip1(\cache_tag[13][21] ), .ip2(addr_resp[29]), .s(n11007), 
        .op(n6984) );
  mux2_1 U11711 ( .ip1(\cache_tag[14][21] ), .ip2(addr_resp[29]), .s(n11008), 
        .op(n6983) );
  mux2_1 U11712 ( .ip1(\cache_tag[15][21] ), .ip2(addr_resp[29]), .s(n11009), 
        .op(n6982) );
  mux2_1 U11713 ( .ip1(N3525), .ip2(addr_req[30]), .s(n7728), .op(n6981) );
  and2_1 U11714 ( .ip1(n11361), .ip2(N3526), .op(n6980) );
  mux2_1 U11715 ( .ip1(\cache_tag[0][22] ), .ip2(addr_resp[30]), .s(n10994), 
        .op(n6979) );
  mux2_1 U11716 ( .ip1(\cache_tag[1][22] ), .ip2(addr_resp[30]), .s(n10995), 
        .op(n6978) );
  mux2_1 U11717 ( .ip1(\cache_tag[2][22] ), .ip2(addr_resp[30]), .s(n10996), 
        .op(n6977) );
  mux2_1 U11718 ( .ip1(\cache_tag[3][22] ), .ip2(addr_resp[30]), .s(n10997), 
        .op(n6976) );
  mux2_1 U11719 ( .ip1(\cache_tag[4][22] ), .ip2(addr_resp[30]), .s(n10998), 
        .op(n6975) );
  mux2_1 U11720 ( .ip1(\cache_tag[5][22] ), .ip2(addr_resp[30]), .s(n10999), 
        .op(n6974) );
  mux2_1 U11721 ( .ip1(\cache_tag[6][22] ), .ip2(addr_resp[30]), .s(n11000), 
        .op(n6973) );
  mux2_1 U11722 ( .ip1(\cache_tag[7][22] ), .ip2(addr_resp[30]), .s(n11001), 
        .op(n6972) );
  mux2_1 U11723 ( .ip1(\cache_tag[8][22] ), .ip2(addr_resp[30]), .s(n11002), 
        .op(n6971) );
  mux2_1 U11724 ( .ip1(\cache_tag[9][22] ), .ip2(addr_resp[30]), .s(n11003), 
        .op(n6970) );
  mux2_1 U11725 ( .ip1(\cache_tag[10][22] ), .ip2(addr_resp[30]), .s(n11004), 
        .op(n6969) );
  mux2_1 U11726 ( .ip1(\cache_tag[11][22] ), .ip2(addr_resp[30]), .s(n11005), 
        .op(n6968) );
  mux2_1 U11727 ( .ip1(\cache_tag[12][22] ), .ip2(addr_resp[30]), .s(n11006), 
        .op(n6967) );
  mux2_1 U11728 ( .ip1(\cache_tag[13][22] ), .ip2(addr_resp[30]), .s(n11007), 
        .op(n6966) );
  mux2_1 U11729 ( .ip1(\cache_tag[14][22] ), .ip2(addr_resp[30]), .s(n11008), 
        .op(n6965) );
  mux2_1 U11730 ( .ip1(\cache_tag[15][22] ), .ip2(addr_resp[30]), .s(n11009), 
        .op(n6964) );
  mux2_1 U11731 ( .ip1(N3522), .ip2(addr_req[31]), .s(n7728), .op(n6963) );
  and2_1 U11732 ( .ip1(n11361), .ip2(N3523), .op(n6962) );
  mux2_1 U11733 ( .ip1(\cache_tag[0][23] ), .ip2(addr_resp[31]), .s(n10994), 
        .op(n6961) );
  mux2_1 U11734 ( .ip1(\cache_tag[1][23] ), .ip2(addr_resp[31]), .s(n10995), 
        .op(n6960) );
  mux2_1 U11735 ( .ip1(\cache_tag[2][23] ), .ip2(addr_resp[31]), .s(n10996), 
        .op(n6959) );
  mux2_1 U11736 ( .ip1(\cache_tag[3][23] ), .ip2(addr_resp[31]), .s(n10997), 
        .op(n6958) );
  mux2_1 U11737 ( .ip1(\cache_tag[4][23] ), .ip2(addr_resp[31]), .s(n10998), 
        .op(n6957) );
  mux2_1 U11738 ( .ip1(\cache_tag[5][23] ), .ip2(addr_resp[31]), .s(n10999), 
        .op(n6956) );
  mux2_1 U11739 ( .ip1(\cache_tag[6][23] ), .ip2(addr_resp[31]), .s(n11000), 
        .op(n6955) );
  mux2_1 U11740 ( .ip1(\cache_tag[7][23] ), .ip2(addr_resp[31]), .s(n11001), 
        .op(n6954) );
  mux2_1 U11741 ( .ip1(\cache_tag[8][23] ), .ip2(addr_resp[31]), .s(n11002), 
        .op(n6953) );
  mux2_1 U11742 ( .ip1(\cache_tag[9][23] ), .ip2(addr_resp[31]), .s(n11003), 
        .op(n6952) );
  mux2_1 U11743 ( .ip1(\cache_tag[10][23] ), .ip2(addr_resp[31]), .s(n11004), 
        .op(n6951) );
  mux2_1 U11744 ( .ip1(\cache_tag[11][23] ), .ip2(addr_resp[31]), .s(n11005), 
        .op(n6950) );
  mux2_1 U11745 ( .ip1(\cache_tag[12][23] ), .ip2(addr_resp[31]), .s(n11006), 
        .op(n6949) );
  mux2_1 U11746 ( .ip1(\cache_tag[13][23] ), .ip2(addr_resp[31]), .s(n11007), 
        .op(n6948) );
  mux2_1 U11747 ( .ip1(\cache_tag[14][23] ), .ip2(addr_resp[31]), .s(n11008), 
        .op(n6947) );
  mux2_1 U11748 ( .ip1(\cache_tag[15][23] ), .ip2(addr_resp[31]), .s(n11009), 
        .op(n6946) );
  nand2_1 U11749 ( .ip1(rd_temp), .ip2(n11361), .op(n11011) );
  nand2_1 U11750 ( .ip1(rd), .ip2(next_state[1]), .op(n11010) );
  nand2_1 U11751 ( .ip1(n11011), .ip2(n11010), .op(n6945) );
  nand2_1 U11752 ( .ip1(rd_temp), .ip2(n12323), .op(n11306) );
  nor3_1 U11753 ( .ip1(addr_resp[2]), .ip2(addr_resp[3]), .ip3(n11306), .op(
        n11293) );
  nand2_1 U11754 ( .ip1(n11293), .ip2(n11012), .op(n11021) );
  inv_1 U11755 ( .ip(addr_resp[2]), .op(n11445) );
  inv_1 U11756 ( .ip(addr_resp[3]), .op(n11444) );
  buf_1 U11757 ( .ip(n11306), .op(n11300) );
  nor3_1 U11758 ( .ip1(n11445), .ip2(n11444), .ip3(n11300), .op(n11302) );
  inv_1 U11759 ( .ip(n11306), .op(n11014) );
  nand3_1 U11760 ( .ip1(addr_resp[3]), .ip2(n11014), .ip3(n11445), .op(n11294)
         );
  nor2_1 U11761 ( .ip1(n11013), .ip2(n11294), .op(n11017) );
  nand3_1 U11762 ( .ip1(addr_resp[2]), .ip2(n11014), .ip3(n11444), .op(n11296)
         );
  nor2_1 U11763 ( .ip1(n11015), .ip2(n11296), .op(n11016) );
  not_ab_or_c_or_d U11764 ( .ip1(n11302), .ip2(n11018), .ip3(n11017), .ip4(
        n11016), .op(n11020) );
  nand2_1 U11765 ( .ip1(N3519), .ip2(n11306), .op(n11019) );
  nand3_1 U11766 ( .ip1(n11021), .ip2(n11020), .ip3(n11019), .op(n6944) );
  and2_1 U11767 ( .ip1(n11306), .ip2(N3520), .op(n6943) );
  nand2_1 U11768 ( .ip1(n11302), .ip2(n11022), .op(n11030) );
  nor2_1 U11769 ( .ip1(n11023), .ip2(n11294), .op(n11026) );
  nor2_1 U11770 ( .ip1(n11024), .ip2(n11296), .op(n11025) );
  not_ab_or_c_or_d U11771 ( .ip1(n11293), .ip2(n11027), .ip3(n11026), .ip4(
        n11025), .op(n11029) );
  nand2_1 U11772 ( .ip1(N3516), .ip2(n11300), .op(n11028) );
  nand3_1 U11773 ( .ip1(n11030), .ip2(n11029), .ip3(n11028), .op(n6942) );
  and2_1 U11774 ( .ip1(n11306), .ip2(N3517), .op(n6941) );
  nand2_1 U11775 ( .ip1(n11293), .ip2(n11031), .op(n11039) );
  nor2_1 U11776 ( .ip1(n11032), .ip2(n11294), .op(n11035) );
  nor2_1 U11777 ( .ip1(n11033), .ip2(n11296), .op(n11034) );
  not_ab_or_c_or_d U11778 ( .ip1(n11302), .ip2(n11036), .ip3(n11035), .ip4(
        n11034), .op(n11038) );
  nand2_1 U11779 ( .ip1(N3513), .ip2(n11306), .op(n11037) );
  nand3_1 U11780 ( .ip1(n11039), .ip2(n11038), .ip3(n11037), .op(n6940) );
  and2_1 U11781 ( .ip1(n11306), .ip2(N3514), .op(n6939) );
  nand2_1 U11782 ( .ip1(n11293), .ip2(n11040), .op(n11048) );
  nor2_1 U11783 ( .ip1(n11041), .ip2(n11296), .op(n11044) );
  nor2_1 U11784 ( .ip1(n11042), .ip2(n11294), .op(n11043) );
  not_ab_or_c_or_d U11785 ( .ip1(n11302), .ip2(n11045), .ip3(n11044), .ip4(
        n11043), .op(n11047) );
  nand2_1 U11786 ( .ip1(N3510), .ip2(n11300), .op(n11046) );
  nand3_1 U11787 ( .ip1(n11048), .ip2(n11047), .ip3(n11046), .op(n6938) );
  and2_1 U11788 ( .ip1(n11306), .ip2(N3511), .op(n6937) );
  nand2_1 U11789 ( .ip1(n11302), .ip2(n11049), .op(n11057) );
  nor2_1 U11790 ( .ip1(n11050), .ip2(n11296), .op(n11053) );
  nor2_1 U11791 ( .ip1(n11051), .ip2(n11294), .op(n11052) );
  not_ab_or_c_or_d U11792 ( .ip1(N3507), .ip2(n11300), .ip3(n11053), .ip4(
        n11052), .op(n11056) );
  nand2_1 U11793 ( .ip1(n11293), .ip2(n11054), .op(n11055) );
  nand3_1 U11794 ( .ip1(n11057), .ip2(n11056), .ip3(n11055), .op(n6936) );
  and2_1 U11795 ( .ip1(n11306), .ip2(N3508), .op(n6935) );
  nand2_1 U11796 ( .ip1(n11302), .ip2(n11058), .op(n11066) );
  nor2_1 U11797 ( .ip1(n11059), .ip2(n11294), .op(n11062) );
  nor2_1 U11798 ( .ip1(n11060), .ip2(n11296), .op(n11061) );
  not_ab_or_c_or_d U11799 ( .ip1(N3504), .ip2(n11300), .ip3(n11062), .ip4(
        n11061), .op(n11065) );
  nand2_1 U11800 ( .ip1(n11293), .ip2(n11063), .op(n11064) );
  nand3_1 U11801 ( .ip1(n11066), .ip2(n11065), .ip3(n11064), .op(n6934) );
  and2_1 U11802 ( .ip1(n11306), .ip2(N3505), .op(n6933) );
  nand2_1 U11803 ( .ip1(n11293), .ip2(n11067), .op(n11075) );
  nor2_1 U11804 ( .ip1(n11068), .ip2(n11294), .op(n11071) );
  nor2_1 U11805 ( .ip1(n11069), .ip2(n11296), .op(n11070) );
  not_ab_or_c_or_d U11806 ( .ip1(n11302), .ip2(n11072), .ip3(n11071), .ip4(
        n11070), .op(n11074) );
  nand2_1 U11807 ( .ip1(N3501), .ip2(n11300), .op(n11073) );
  nand3_1 U11808 ( .ip1(n11075), .ip2(n11074), .ip3(n11073), .op(n6932) );
  and2_1 U11809 ( .ip1(n11306), .ip2(N3502), .op(n6931) );
  nand2_1 U11810 ( .ip1(n11293), .ip2(n11076), .op(n11084) );
  nor2_1 U11811 ( .ip1(n11077), .ip2(n11294), .op(n11080) );
  nor2_1 U11812 ( .ip1(n11078), .ip2(n11296), .op(n11079) );
  not_ab_or_c_or_d U11813 ( .ip1(n11302), .ip2(n11081), .ip3(n11080), .ip4(
        n11079), .op(n11083) );
  nand2_1 U11814 ( .ip1(N3498), .ip2(n11300), .op(n11082) );
  nand3_1 U11815 ( .ip1(n11084), .ip2(n11083), .ip3(n11082), .op(n6930) );
  and2_1 U11816 ( .ip1(n11306), .ip2(N3499), .op(n6929) );
  nand2_1 U11817 ( .ip1(n11293), .ip2(n11085), .op(n11093) );
  nor2_1 U11818 ( .ip1(n11086), .ip2(n11294), .op(n11089) );
  nor2_1 U11819 ( .ip1(n11087), .ip2(n11296), .op(n11088) );
  not_ab_or_c_or_d U11820 ( .ip1(N3495), .ip2(n11300), .ip3(n11089), .ip4(
        n11088), .op(n11092) );
  nand2_1 U11821 ( .ip1(n11302), .ip2(n11090), .op(n11091) );
  nand3_1 U11822 ( .ip1(n11093), .ip2(n11092), .ip3(n11091), .op(n6928) );
  and2_1 U11823 ( .ip1(n11306), .ip2(N3496), .op(n6927) );
  nand2_1 U11824 ( .ip1(n11302), .ip2(n11094), .op(n11102) );
  nor2_1 U11825 ( .ip1(n11095), .ip2(n11294), .op(n11098) );
  nor2_1 U11826 ( .ip1(n11096), .ip2(n11296), .op(n11097) );
  not_ab_or_c_or_d U11827 ( .ip1(n11293), .ip2(n11099), .ip3(n11098), .ip4(
        n11097), .op(n11101) );
  nand2_1 U11828 ( .ip1(N3492), .ip2(n11306), .op(n11100) );
  nand3_1 U11829 ( .ip1(n11102), .ip2(n11101), .ip3(n11100), .op(n6926) );
  and2_1 U11830 ( .ip1(n11306), .ip2(N3493), .op(n6925) );
  nand2_1 U11831 ( .ip1(n11293), .ip2(n11103), .op(n11111) );
  nor2_1 U11832 ( .ip1(n11104), .ip2(n11294), .op(n11107) );
  nor2_1 U11833 ( .ip1(n11105), .ip2(n11296), .op(n11106) );
  not_ab_or_c_or_d U11834 ( .ip1(N3489), .ip2(n11300), .ip3(n11107), .ip4(
        n11106), .op(n11110) );
  nand2_1 U11835 ( .ip1(n11302), .ip2(n11108), .op(n11109) );
  nand3_1 U11836 ( .ip1(n11111), .ip2(n11110), .ip3(n11109), .op(n6924) );
  and2_1 U11837 ( .ip1(n11306), .ip2(N3490), .op(n6923) );
  nand2_1 U11838 ( .ip1(n11293), .ip2(n11112), .op(n11120) );
  nor2_1 U11839 ( .ip1(n11113), .ip2(n11296), .op(n11116) );
  nor2_1 U11840 ( .ip1(n11114), .ip2(n11294), .op(n11115) );
  not_ab_or_c_or_d U11841 ( .ip1(n11302), .ip2(n11117), .ip3(n11116), .ip4(
        n11115), .op(n11119) );
  nand2_1 U11842 ( .ip1(N3486), .ip2(n11300), .op(n11118) );
  nand3_1 U11843 ( .ip1(n11120), .ip2(n11119), .ip3(n11118), .op(n6922) );
  and2_1 U11844 ( .ip1(n11306), .ip2(N3487), .op(n6921) );
  nand2_1 U11845 ( .ip1(n11302), .ip2(n11121), .op(n11129) );
  nor2_1 U11846 ( .ip1(n11122), .ip2(n11294), .op(n11125) );
  nor2_1 U11847 ( .ip1(n11123), .ip2(n11296), .op(n11124) );
  not_ab_or_c_or_d U11848 ( .ip1(N3483), .ip2(n11300), .ip3(n11125), .ip4(
        n11124), .op(n11128) );
  nand2_1 U11849 ( .ip1(n11293), .ip2(n11126), .op(n11127) );
  nand3_1 U11850 ( .ip1(n11129), .ip2(n11128), .ip3(n11127), .op(n6920) );
  and2_1 U11851 ( .ip1(n11306), .ip2(N3484), .op(n6919) );
  nand2_1 U11852 ( .ip1(n11293), .ip2(n11130), .op(n11138) );
  nor2_1 U11853 ( .ip1(n11131), .ip2(n11294), .op(n11134) );
  nor2_1 U11854 ( .ip1(n11132), .ip2(n11296), .op(n11133) );
  not_ab_or_c_or_d U11855 ( .ip1(n11302), .ip2(n11135), .ip3(n11134), .ip4(
        n11133), .op(n11137) );
  nand2_1 U11856 ( .ip1(N3480), .ip2(n11300), .op(n11136) );
  nand3_1 U11857 ( .ip1(n11138), .ip2(n11137), .ip3(n11136), .op(n6918) );
  and2_1 U11858 ( .ip1(n11306), .ip2(N3481), .op(n6917) );
  nand2_1 U11859 ( .ip1(n11293), .ip2(n11139), .op(n11147) );
  nor2_1 U11860 ( .ip1(n11140), .ip2(n11296), .op(n11143) );
  nor2_1 U11861 ( .ip1(n11141), .ip2(n11294), .op(n11142) );
  not_ab_or_c_or_d U11862 ( .ip1(n11302), .ip2(n11144), .ip3(n11143), .ip4(
        n11142), .op(n11146) );
  nand2_1 U11863 ( .ip1(N3477), .ip2(n11300), .op(n11145) );
  nand3_1 U11864 ( .ip1(n11147), .ip2(n11146), .ip3(n11145), .op(n6916) );
  and2_1 U11865 ( .ip1(n11306), .ip2(N3478), .op(n6915) );
  nand2_1 U11866 ( .ip1(n11293), .ip2(n11148), .op(n11156) );
  nor2_1 U11867 ( .ip1(n11149), .ip2(n11294), .op(n11152) );
  nor2_1 U11868 ( .ip1(n11150), .ip2(n11296), .op(n11151) );
  not_ab_or_c_or_d U11869 ( .ip1(n11302), .ip2(n11153), .ip3(n11152), .ip4(
        n11151), .op(n11155) );
  nand2_1 U11870 ( .ip1(N3474), .ip2(n11300), .op(n11154) );
  nand3_1 U11871 ( .ip1(n11156), .ip2(n11155), .ip3(n11154), .op(n6914) );
  and2_1 U11872 ( .ip1(n11306), .ip2(N3475), .op(n6913) );
  nand2_1 U11873 ( .ip1(n11293), .ip2(n11157), .op(n11165) );
  nor2_1 U11874 ( .ip1(n11158), .ip2(n11294), .op(n11161) );
  nor2_1 U11875 ( .ip1(n11159), .ip2(n11296), .op(n11160) );
  not_ab_or_c_or_d U11876 ( .ip1(n11302), .ip2(n11162), .ip3(n11161), .ip4(
        n11160), .op(n11164) );
  nand2_1 U11877 ( .ip1(N3471), .ip2(n11300), .op(n11163) );
  nand3_1 U11878 ( .ip1(n11165), .ip2(n11164), .ip3(n11163), .op(n6912) );
  and2_1 U11879 ( .ip1(n11306), .ip2(N3472), .op(n6911) );
  nand2_1 U11880 ( .ip1(n11302), .ip2(n11166), .op(n11174) );
  nor2_1 U11881 ( .ip1(n11167), .ip2(n11296), .op(n11170) );
  nor2_1 U11882 ( .ip1(n11168), .ip2(n11294), .op(n11169) );
  not_ab_or_c_or_d U11883 ( .ip1(N3468), .ip2(n11300), .ip3(n11170), .ip4(
        n11169), .op(n11173) );
  nand2_1 U11884 ( .ip1(n11293), .ip2(n11171), .op(n11172) );
  nand3_1 U11885 ( .ip1(n11174), .ip2(n11173), .ip3(n11172), .op(n6910) );
  and2_1 U11886 ( .ip1(n11306), .ip2(N3469), .op(n6909) );
  nand2_1 U11887 ( .ip1(n11293), .ip2(n11175), .op(n11183) );
  nor2_1 U11888 ( .ip1(n11176), .ip2(n11296), .op(n11179) );
  nor2_1 U11889 ( .ip1(n11177), .ip2(n11294), .op(n11178) );
  not_ab_or_c_or_d U11890 ( .ip1(n11302), .ip2(n11180), .ip3(n11179), .ip4(
        n11178), .op(n11182) );
  nand2_1 U11891 ( .ip1(N3465), .ip2(n11306), .op(n11181) );
  nand3_1 U11892 ( .ip1(n11183), .ip2(n11182), .ip3(n11181), .op(n6908) );
  and2_1 U11893 ( .ip1(n11306), .ip2(N3466), .op(n6907) );
  nand2_1 U11894 ( .ip1(n11293), .ip2(n11184), .op(n11192) );
  nor2_1 U11895 ( .ip1(n11185), .ip2(n11294), .op(n11188) );
  nor2_1 U11896 ( .ip1(n11186), .ip2(n11296), .op(n11187) );
  not_ab_or_c_or_d U11897 ( .ip1(N3462), .ip2(n11300), .ip3(n11188), .ip4(
        n11187), .op(n11191) );
  nand2_1 U11898 ( .ip1(n11302), .ip2(n11189), .op(n11190) );
  nand3_1 U11899 ( .ip1(n11192), .ip2(n11191), .ip3(n11190), .op(n6906) );
  and2_1 U11900 ( .ip1(n11306), .ip2(N3463), .op(n6905) );
  nand2_1 U11901 ( .ip1(n11293), .ip2(n11193), .op(n11201) );
  nor2_1 U11902 ( .ip1(n11194), .ip2(n11296), .op(n11197) );
  nor2_1 U11903 ( .ip1(n11195), .ip2(n11294), .op(n11196) );
  not_ab_or_c_or_d U11904 ( .ip1(N3459), .ip2(n11300), .ip3(n11197), .ip4(
        n11196), .op(n11200) );
  nand2_1 U11905 ( .ip1(n11302), .ip2(n11198), .op(n11199) );
  nand3_1 U11906 ( .ip1(n11201), .ip2(n11200), .ip3(n11199), .op(n6904) );
  and2_1 U11907 ( .ip1(n11306), .ip2(N3460), .op(n6903) );
  nand2_1 U11908 ( .ip1(n11302), .ip2(n11202), .op(n11210) );
  nor2_1 U11909 ( .ip1(n11203), .ip2(n11296), .op(n11206) );
  nor2_1 U11910 ( .ip1(n11204), .ip2(n11294), .op(n11205) );
  not_ab_or_c_or_d U11911 ( .ip1(n11293), .ip2(n11207), .ip3(n11206), .ip4(
        n11205), .op(n11209) );
  nand2_1 U11912 ( .ip1(N3456), .ip2(n11306), .op(n11208) );
  nand3_1 U11913 ( .ip1(n11210), .ip2(n11209), .ip3(n11208), .op(n6902) );
  and2_1 U11914 ( .ip1(n11306), .ip2(N3457), .op(n6901) );
  nand2_1 U11915 ( .ip1(n11302), .ip2(n11211), .op(n11219) );
  nor2_1 U11916 ( .ip1(n11212), .ip2(n11294), .op(n11215) );
  nor2_1 U11917 ( .ip1(n11213), .ip2(n11296), .op(n11214) );
  not_ab_or_c_or_d U11918 ( .ip1(N3453), .ip2(n11300), .ip3(n11215), .ip4(
        n11214), .op(n11218) );
  nand2_1 U11919 ( .ip1(n11293), .ip2(n11216), .op(n11217) );
  nand3_1 U11920 ( .ip1(n11219), .ip2(n11218), .ip3(n11217), .op(n6900) );
  and2_1 U11921 ( .ip1(n11306), .ip2(N3454), .op(n6899) );
  nand2_1 U11922 ( .ip1(n11302), .ip2(n11220), .op(n11228) );
  nor2_1 U11923 ( .ip1(n11221), .ip2(n11294), .op(n11224) );
  nor2_1 U11924 ( .ip1(n11222), .ip2(n11296), .op(n11223) );
  not_ab_or_c_or_d U11925 ( .ip1(n11293), .ip2(n11225), .ip3(n11224), .ip4(
        n11223), .op(n11227) );
  nand2_1 U11926 ( .ip1(N3450), .ip2(n11306), .op(n11226) );
  nand3_1 U11927 ( .ip1(n11228), .ip2(n11227), .ip3(n11226), .op(n6898) );
  and2_1 U11928 ( .ip1(n11306), .ip2(N3451), .op(n6897) );
  nand2_1 U11929 ( .ip1(n11293), .ip2(n11229), .op(n11237) );
  nor2_1 U11930 ( .ip1(n11230), .ip2(n11294), .op(n11233) );
  nor2_1 U11931 ( .ip1(n11231), .ip2(n11296), .op(n11232) );
  not_ab_or_c_or_d U11932 ( .ip1(n11302), .ip2(n11234), .ip3(n11233), .ip4(
        n11232), .op(n11236) );
  nand2_1 U11933 ( .ip1(N3447), .ip2(n11306), .op(n11235) );
  nand3_1 U11934 ( .ip1(n11237), .ip2(n11236), .ip3(n11235), .op(n6896) );
  and2_1 U11935 ( .ip1(n11306), .ip2(N3448), .op(n6895) );
  nand2_1 U11936 ( .ip1(n11302), .ip2(n11238), .op(n11246) );
  nor2_1 U11937 ( .ip1(n11239), .ip2(n11294), .op(n11242) );
  nor2_1 U11938 ( .ip1(n11240), .ip2(n11296), .op(n11241) );
  not_ab_or_c_or_d U11939 ( .ip1(N3444), .ip2(n11300), .ip3(n11242), .ip4(
        n11241), .op(n11245) );
  nand2_1 U11940 ( .ip1(n11293), .ip2(n11243), .op(n11244) );
  nand3_1 U11941 ( .ip1(n11246), .ip2(n11245), .ip3(n11244), .op(n6894) );
  and2_1 U11942 ( .ip1(n11306), .ip2(N3445), .op(n6893) );
  nand2_1 U11943 ( .ip1(n11302), .ip2(n11247), .op(n11255) );
  nor2_1 U11944 ( .ip1(n11248), .ip2(n11296), .op(n11251) );
  nor2_1 U11945 ( .ip1(n11249), .ip2(n11294), .op(n11250) );
  not_ab_or_c_or_d U11946 ( .ip1(N3441), .ip2(n11300), .ip3(n11251), .ip4(
        n11250), .op(n11254) );
  nand2_1 U11947 ( .ip1(n11293), .ip2(n11252), .op(n11253) );
  nand3_1 U11948 ( .ip1(n11255), .ip2(n11254), .ip3(n11253), .op(n6892) );
  and2_1 U11949 ( .ip1(n11306), .ip2(N3442), .op(n6891) );
  nand2_1 U11950 ( .ip1(n11302), .ip2(n11256), .op(n11264) );
  nor2_1 U11951 ( .ip1(n11257), .ip2(n11296), .op(n11260) );
  nor2_1 U11952 ( .ip1(n11258), .ip2(n11294), .op(n11259) );
  not_ab_or_c_or_d U11953 ( .ip1(N3438), .ip2(n11300), .ip3(n11260), .ip4(
        n11259), .op(n11263) );
  nand2_1 U11954 ( .ip1(n11293), .ip2(n11261), .op(n11262) );
  nand3_1 U11955 ( .ip1(n11264), .ip2(n11263), .ip3(n11262), .op(n6890) );
  and2_1 U11956 ( .ip1(n11306), .ip2(N3439), .op(n6889) );
  nand2_1 U11957 ( .ip1(n11302), .ip2(n11265), .op(n11273) );
  nor2_1 U11958 ( .ip1(n11266), .ip2(n11296), .op(n11269) );
  nor2_1 U11959 ( .ip1(n11267), .ip2(n11294), .op(n11268) );
  not_ab_or_c_or_d U11960 ( .ip1(N3435), .ip2(n11300), .ip3(n11269), .ip4(
        n11268), .op(n11272) );
  nand2_1 U11961 ( .ip1(n11293), .ip2(n11270), .op(n11271) );
  nand3_1 U11962 ( .ip1(n11273), .ip2(n11272), .ip3(n11271), .op(n6888) );
  and2_1 U11963 ( .ip1(n11306), .ip2(N3436), .op(n6887) );
  nand2_1 U11964 ( .ip1(n11302), .ip2(n11274), .op(n11282) );
  nor2_1 U11965 ( .ip1(n11275), .ip2(n11296), .op(n11278) );
  nor2_1 U11966 ( .ip1(n11276), .ip2(n11294), .op(n11277) );
  not_ab_or_c_or_d U11967 ( .ip1(n11293), .ip2(n11279), .ip3(n11278), .ip4(
        n11277), .op(n11281) );
  nand2_1 U11968 ( .ip1(N3432), .ip2(n11306), .op(n11280) );
  nand3_1 U11969 ( .ip1(n11282), .ip2(n11281), .ip3(n11280), .op(n6886) );
  and2_1 U11970 ( .ip1(n11306), .ip2(N3433), .op(n6885) );
  nand2_1 U11971 ( .ip1(n11293), .ip2(n11283), .op(n11291) );
  nor2_1 U11972 ( .ip1(n11284), .ip2(n11296), .op(n11287) );
  nor2_1 U11973 ( .ip1(n11285), .ip2(n11294), .op(n11286) );
  not_ab_or_c_or_d U11974 ( .ip1(N3429), .ip2(n11300), .ip3(n11287), .ip4(
        n11286), .op(n11290) );
  nand2_1 U11975 ( .ip1(n11302), .ip2(n11288), .op(n11289) );
  nand3_1 U11976 ( .ip1(n11291), .ip2(n11290), .ip3(n11289), .op(n6884) );
  and2_1 U11977 ( .ip1(n11306), .ip2(N3430), .op(n6883) );
  nand2_1 U11978 ( .ip1(n11293), .ip2(n11292), .op(n11305) );
  nor2_1 U11979 ( .ip1(n11295), .ip2(n11294), .op(n11299) );
  nor2_1 U11980 ( .ip1(n11297), .ip2(n11296), .op(n11298) );
  not_ab_or_c_or_d U11981 ( .ip1(N3426), .ip2(n11300), .ip3(n11299), .ip4(
        n11298), .op(n11304) );
  nand2_1 U11982 ( .ip1(n11302), .ip2(n11301), .op(n11303) );
  nand3_1 U11983 ( .ip1(n11305), .ip2(n11304), .ip3(n11303), .op(n6882) );
  and2_1 U11984 ( .ip1(n11306), .ip2(N3427), .op(n6881) );
  nor2_1 U11985 ( .ip1(n11307), .ip2(rd_temp), .op(n11366) );
  nand2_1 U11986 ( .ip1(n11964), .ip2(n11366), .op(n11310) );
  nand2_1 U11987 ( .ip1(cache_dirty[0]), .ip2(n11308), .op(n11309) );
  nand2_1 U11988 ( .ip1(n11310), .ip2(n11309), .op(n6880) );
  nand2_1 U11989 ( .ip1(n11943), .ip2(n11366), .op(n11313) );
  nand2_1 U11990 ( .ip1(cache_dirty[1]), .ip2(n11311), .op(n11312) );
  nand2_1 U11991 ( .ip1(n11313), .ip2(n11312), .op(n6879) );
  nand2_1 U11992 ( .ip1(n12228), .ip2(n11366), .op(n11316) );
  nand2_1 U11993 ( .ip1(cache_dirty[2]), .ip2(n11314), .op(n11315) );
  nand2_1 U11994 ( .ip1(n11316), .ip2(n11315), .op(n6878) );
  nand2_1 U11995 ( .ip1(n11317), .ip2(n11366), .op(n11320) );
  nand2_1 U11996 ( .ip1(cache_dirty[3]), .ip2(n11318), .op(n11319) );
  nand2_1 U11997 ( .ip1(n11320), .ip2(n11319), .op(n6877) );
  nand2_1 U11998 ( .ip1(n12164), .ip2(n11366), .op(n11323) );
  nand2_1 U11999 ( .ip1(cache_dirty[4]), .ip2(n11321), .op(n11322) );
  nand2_1 U12000 ( .ip1(n11323), .ip2(n11322), .op(n6876) );
  nand2_1 U12001 ( .ip1(n11963), .ip2(n11366), .op(n11326) );
  nand2_1 U12002 ( .ip1(cache_dirty[5]), .ip2(n11324), .op(n11325) );
  nand2_1 U12003 ( .ip1(n11326), .ip2(n11325), .op(n6875) );
  nand2_1 U12004 ( .ip1(n11972), .ip2(n11366), .op(n11329) );
  nand2_1 U12005 ( .ip1(cache_dirty[6]), .ip2(n11327), .op(n11328) );
  nand2_1 U12006 ( .ip1(n11329), .ip2(n11328), .op(n6874) );
  nand2_1 U12007 ( .ip1(n12202), .ip2(n11366), .op(n11332) );
  nand2_1 U12008 ( .ip1(cache_dirty[7]), .ip2(n11330), .op(n11331) );
  nand2_1 U12009 ( .ip1(n11332), .ip2(n11331), .op(n6873) );
  nand2_1 U12010 ( .ip1(n12234), .ip2(n11366), .op(n11335) );
  nand2_1 U12011 ( .ip1(cache_dirty[8]), .ip2(n11333), .op(n11334) );
  nand2_1 U12012 ( .ip1(n11335), .ip2(n11334), .op(n6872) );
  nand2_1 U12013 ( .ip1(n12241), .ip2(n11366), .op(n11338) );
  nand2_1 U12014 ( .ip1(cache_dirty[9]), .ip2(n11336), .op(n11337) );
  nand2_1 U12015 ( .ip1(n11338), .ip2(n11337), .op(n6871) );
  nand2_1 U12016 ( .ip1(n11966), .ip2(n11366), .op(n11341) );
  nand2_1 U12017 ( .ip1(cache_dirty[10]), .ip2(n11339), .op(n11340) );
  nand2_1 U12018 ( .ip1(n11341), .ip2(n11340), .op(n6870) );
  nand2_1 U12019 ( .ip1(n12170), .ip2(n11366), .op(n11344) );
  nand2_1 U12020 ( .ip1(cache_dirty[11]), .ip2(n11342), .op(n11343) );
  nand2_1 U12021 ( .ip1(n11344), .ip2(n11343), .op(n6869) );
  nand2_1 U12022 ( .ip1(n12030), .ip2(n11366), .op(n11347) );
  nand2_1 U12023 ( .ip1(cache_dirty[12]), .ip2(n11345), .op(n11346) );
  nand2_1 U12024 ( .ip1(n11347), .ip2(n11346), .op(n6868) );
  nand2_1 U12025 ( .ip1(n12242), .ip2(n11366), .op(n11350) );
  nand2_1 U12026 ( .ip1(cache_dirty[13]), .ip2(n11348), .op(n11349) );
  nand2_1 U12027 ( .ip1(n11350), .ip2(n11349), .op(n6867) );
  nand2_1 U12028 ( .ip1(n11688), .ip2(n11366), .op(n11353) );
  nand2_1 U12029 ( .ip1(cache_dirty[14]), .ip2(n11351), .op(n11352) );
  nand2_1 U12030 ( .ip1(n11353), .ip2(n11352), .op(n6866) );
  nand2_1 U12031 ( .ip1(n11965), .ip2(n11366), .op(n11356) );
  nand2_1 U12032 ( .ip1(cache_dirty[15]), .ip2(n11354), .op(n11355) );
  nand2_1 U12033 ( .ip1(n11356), .ip2(n11355), .op(n6865) );
  nor2_1 U12034 ( .ip1(n11358), .ip2(n11357), .op(n11359) );
  or2_1 U12035 ( .ip1(n11360), .ip2(n11359), .op(n6864) );
  nor2_1 U12036 ( .ip1(rst), .ip2(n11361), .op(n11362) );
  buf_1 U12037 ( .ip(n11362), .op(n11363) );
  mux2_1 U12038 ( .ip1(iCache_data_wr[0]), .ip2(data_wr[0]), .s(n11363), .op(
        n6863) );
  mux2_1 U12039 ( .ip1(iCache_data_wr[1]), .ip2(data_wr[1]), .s(n11362), .op(
        n6862) );
  mux2_1 U12040 ( .ip1(iCache_data_wr[2]), .ip2(data_wr[2]), .s(n11362), .op(
        n6861) );
  mux2_1 U12041 ( .ip1(iCache_data_wr[3]), .ip2(data_wr[3]), .s(n11362), .op(
        n6860) );
  mux2_1 U12042 ( .ip1(iCache_data_wr[4]), .ip2(data_wr[4]), .s(n11362), .op(
        n6859) );
  mux2_1 U12043 ( .ip1(iCache_data_wr[5]), .ip2(data_wr[5]), .s(n11362), .op(
        n6858) );
  mux2_1 U12044 ( .ip1(iCache_data_wr[6]), .ip2(data_wr[6]), .s(n11362), .op(
        n6857) );
  mux2_1 U12045 ( .ip1(iCache_data_wr[7]), .ip2(data_wr[7]), .s(n11362), .op(
        n6856) );
  mux2_1 U12046 ( .ip1(iCache_data_wr[8]), .ip2(data_wr[8]), .s(n11362), .op(
        n6855) );
  mux2_1 U12047 ( .ip1(iCache_data_wr[9]), .ip2(data_wr[9]), .s(n11363), .op(
        n6854) );
  mux2_1 U12048 ( .ip1(iCache_data_wr[10]), .ip2(data_wr[10]), .s(n11363), 
        .op(n6853) );
  mux2_1 U12049 ( .ip1(iCache_data_wr[11]), .ip2(data_wr[11]), .s(n11362), 
        .op(n6852) );
  mux2_1 U12050 ( .ip1(iCache_data_wr[12]), .ip2(data_wr[12]), .s(n11362), 
        .op(n6851) );
  mux2_1 U12051 ( .ip1(iCache_data_wr[13]), .ip2(data_wr[13]), .s(n11362), 
        .op(n6850) );
  mux2_1 U12052 ( .ip1(iCache_data_wr[14]), .ip2(data_wr[14]), .s(n11362), 
        .op(n6849) );
  mux2_1 U12053 ( .ip1(iCache_data_wr[15]), .ip2(data_wr[15]), .s(n11362), 
        .op(n6848) );
  mux2_1 U12054 ( .ip1(iCache_data_wr[16]), .ip2(data_wr[16]), .s(n11362), 
        .op(n6847) );
  mux2_1 U12055 ( .ip1(iCache_data_wr[17]), .ip2(data_wr[17]), .s(n11362), 
        .op(n6846) );
  mux2_1 U12056 ( .ip1(iCache_data_wr[18]), .ip2(data_wr[18]), .s(n11362), 
        .op(n6845) );
  mux2_1 U12057 ( .ip1(iCache_data_wr[19]), .ip2(data_wr[19]), .s(n11362), 
        .op(n6844) );
  mux2_1 U12058 ( .ip1(iCache_data_wr[20]), .ip2(data_wr[20]), .s(n11362), 
        .op(n6843) );
  mux2_1 U12059 ( .ip1(iCache_data_wr[21]), .ip2(data_wr[21]), .s(n11362), 
        .op(n6842) );
  mux2_1 U12060 ( .ip1(iCache_data_wr[22]), .ip2(data_wr[22]), .s(n11362), 
        .op(n6841) );
  mux2_1 U12061 ( .ip1(iCache_data_wr[23]), .ip2(data_wr[23]), .s(n11362), 
        .op(n6840) );
  mux2_1 U12062 ( .ip1(iCache_data_wr[24]), .ip2(data_wr[24]), .s(n11363), 
        .op(n6839) );
  mux2_1 U12063 ( .ip1(iCache_data_wr[25]), .ip2(data_wr[25]), .s(n11363), 
        .op(n6838) );
  mux2_1 U12064 ( .ip1(iCache_data_wr[26]), .ip2(data_wr[26]), .s(n11363), 
        .op(n6837) );
  mux2_1 U12065 ( .ip1(iCache_data_wr[27]), .ip2(data_wr[27]), .s(n11363), 
        .op(n6836) );
  mux2_1 U12066 ( .ip1(iCache_data_wr[28]), .ip2(data_wr[28]), .s(n11363), 
        .op(n6835) );
  mux2_1 U12067 ( .ip1(iCache_data_wr[29]), .ip2(data_wr[29]), .s(n11363), 
        .op(n6834) );
  mux2_1 U12068 ( .ip1(iCache_data_wr[30]), .ip2(data_wr[30]), .s(n11363), 
        .op(n6833) );
  mux2_1 U12069 ( .ip1(iCache_data_wr[31]), .ip2(data_wr[31]), .s(n11363), 
        .op(n6832) );
  nand2_1 U12070 ( .ip1(iCache_data_wr[0]), .ip2(n12323), .op(n11365) );
  nand2_1 U12071 ( .ip1(data_rd_mem[0]), .ip2(n12325), .op(n11364) );
  nand2_1 U12072 ( .ip1(n11365), .ip2(n11364), .op(n11554) );
  nand2_1 U12073 ( .ip1(n11366), .ip2(n12326), .op(n11446) );
  nor3_1 U12074 ( .ip1(addr_resp[2]), .ip2(addr_resp[3]), .ip3(n11446), .op(
        n11368) );
  nand2_1 U12075 ( .ip1(n12254), .ip2(n12326), .op(n11443) );
  nor3_1 U12076 ( .ip1(mem_data_cnt[2]), .ip2(n11443), .ip3(mem_data_cnt[3]), 
        .op(n11367) );
  nor2_1 U12077 ( .ip1(n11368), .ip2(n11367), .op(n11603) );
  nor2_1 U12078 ( .ip1(n11603), .ip2(n8923), .op(n11415) );
  mux2_1 U12079 ( .ip1(\cache_data[0][0] ), .ip2(n11554), .s(n11415), .op(
        n6831) );
  nand2_1 U12080 ( .ip1(iCache_data_wr[1]), .ip2(n12323), .op(n11370) );
  nand2_1 U12081 ( .ip1(data_rd_mem[1]), .ip2(n12325), .op(n11369) );
  nand2_1 U12082 ( .ip1(n11370), .ip2(n11369), .op(n11555) );
  mux2_1 U12083 ( .ip1(\cache_data[0][1] ), .ip2(n11555), .s(n11415), .op(
        n6830) );
  nand2_1 U12084 ( .ip1(iCache_data_wr[2]), .ip2(n12323), .op(n11372) );
  nand2_1 U12085 ( .ip1(data_rd_mem[2]), .ip2(n12325), .op(n11371) );
  nand2_1 U12086 ( .ip1(n11372), .ip2(n11371), .op(n11556) );
  mux2_1 U12087 ( .ip1(\cache_data[0][2] ), .ip2(n11556), .s(n11415), .op(
        n6829) );
  nand2_1 U12088 ( .ip1(iCache_data_wr[3]), .ip2(n12323), .op(n11374) );
  nand2_1 U12089 ( .ip1(data_rd_mem[3]), .ip2(n12325), .op(n11373) );
  nand2_1 U12090 ( .ip1(n11374), .ip2(n11373), .op(n11557) );
  mux2_1 U12091 ( .ip1(\cache_data[0][3] ), .ip2(n11557), .s(n11415), .op(
        n6828) );
  nand2_1 U12092 ( .ip1(iCache_data_wr[4]), .ip2(n12323), .op(n11376) );
  nand2_1 U12093 ( .ip1(data_rd_mem[4]), .ip2(n12325), .op(n11375) );
  nand2_1 U12094 ( .ip1(n11376), .ip2(n11375), .op(n11558) );
  mux2_1 U12095 ( .ip1(\cache_data[0][4] ), .ip2(n11558), .s(n11415), .op(
        n6827) );
  nand2_1 U12096 ( .ip1(iCache_data_wr[5]), .ip2(n12323), .op(n11378) );
  nand2_1 U12097 ( .ip1(data_rd_mem[5]), .ip2(n12325), .op(n11377) );
  nand2_1 U12098 ( .ip1(n11378), .ip2(n11377), .op(n11559) );
  mux2_1 U12099 ( .ip1(\cache_data[0][5] ), .ip2(n11559), .s(n11415), .op(
        n6826) );
  nand2_1 U12100 ( .ip1(iCache_data_wr[6]), .ip2(n12323), .op(n11380) );
  nand2_1 U12101 ( .ip1(data_rd_mem[6]), .ip2(n12325), .op(n11379) );
  nand2_1 U12102 ( .ip1(n11380), .ip2(n11379), .op(n11560) );
  mux2_1 U12103 ( .ip1(\cache_data[0][6] ), .ip2(n11560), .s(n11415), .op(
        n6825) );
  nand2_1 U12104 ( .ip1(iCache_data_wr[7]), .ip2(n12323), .op(n11382) );
  nand2_1 U12105 ( .ip1(data_rd_mem[7]), .ip2(n12325), .op(n11381) );
  nand2_1 U12106 ( .ip1(n11382), .ip2(n11381), .op(n11561) );
  mux2_1 U12107 ( .ip1(\cache_data[0][7] ), .ip2(n11561), .s(n11415), .op(
        n6824) );
  nand2_1 U12108 ( .ip1(iCache_data_wr[8]), .ip2(n12323), .op(n11384) );
  nand2_1 U12109 ( .ip1(data_rd_mem[8]), .ip2(n12325), .op(n11383) );
  nand2_1 U12110 ( .ip1(n11384), .ip2(n11383), .op(n11562) );
  mux2_1 U12111 ( .ip1(\cache_data[0][8] ), .ip2(n11562), .s(n11415), .op(
        n6823) );
  nand2_1 U12112 ( .ip1(iCache_data_wr[9]), .ip2(n12323), .op(n11386) );
  nand2_1 U12113 ( .ip1(data_rd_mem[9]), .ip2(n12325), .op(n11385) );
  nand2_1 U12114 ( .ip1(n11386), .ip2(n11385), .op(n11563) );
  buf_1 U12115 ( .ip(n11415), .op(n11432) );
  mux2_1 U12116 ( .ip1(\cache_data[0][9] ), .ip2(n11563), .s(n11432), .op(
        n6822) );
  nand2_1 U12117 ( .ip1(iCache_data_wr[10]), .ip2(n12323), .op(n11388) );
  nand2_1 U12118 ( .ip1(data_rd_mem[10]), .ip2(n12325), .op(n11387) );
  nand2_1 U12119 ( .ip1(n11388), .ip2(n11387), .op(n11564) );
  mux2_1 U12120 ( .ip1(\cache_data[0][10] ), .ip2(n11564), .s(n11432), .op(
        n6821) );
  nand2_1 U12121 ( .ip1(iCache_data_wr[11]), .ip2(n12323), .op(n11390) );
  nand2_1 U12122 ( .ip1(data_rd_mem[11]), .ip2(n12325), .op(n11389) );
  nand2_1 U12123 ( .ip1(n11390), .ip2(n11389), .op(n11565) );
  mux2_1 U12124 ( .ip1(\cache_data[0][11] ), .ip2(n11565), .s(n11415), .op(
        n6820) );
  nand2_1 U12125 ( .ip1(iCache_data_wr[12]), .ip2(n12323), .op(n11392) );
  nand2_1 U12126 ( .ip1(data_rd_mem[12]), .ip2(n12325), .op(n11391) );
  nand2_1 U12127 ( .ip1(n11392), .ip2(n11391), .op(n11566) );
  mux2_1 U12128 ( .ip1(\cache_data[0][12] ), .ip2(n11566), .s(n11415), .op(
        n6819) );
  nand2_1 U12129 ( .ip1(iCache_data_wr[13]), .ip2(n12323), .op(n11394) );
  nand2_1 U12130 ( .ip1(data_rd_mem[13]), .ip2(n12325), .op(n11393) );
  nand2_1 U12131 ( .ip1(n11394), .ip2(n11393), .op(n11567) );
  mux2_1 U12132 ( .ip1(\cache_data[0][13] ), .ip2(n11567), .s(n11432), .op(
        n6818) );
  nand2_1 U12133 ( .ip1(iCache_data_wr[14]), .ip2(n12323), .op(n11396) );
  nand2_1 U12134 ( .ip1(data_rd_mem[14]), .ip2(n12325), .op(n11395) );
  nand2_1 U12135 ( .ip1(n11396), .ip2(n11395), .op(n11568) );
  mux2_1 U12136 ( .ip1(\cache_data[0][14] ), .ip2(n11568), .s(n11415), .op(
        n6817) );
  nand2_1 U12137 ( .ip1(iCache_data_wr[15]), .ip2(n12323), .op(n11398) );
  nand2_1 U12138 ( .ip1(data_rd_mem[15]), .ip2(n12325), .op(n11397) );
  nand2_1 U12139 ( .ip1(n11398), .ip2(n11397), .op(n11569) );
  mux2_1 U12140 ( .ip1(\cache_data[0][15] ), .ip2(n11569), .s(n11415), .op(
        n6816) );
  nand2_1 U12141 ( .ip1(iCache_data_wr[16]), .ip2(n12323), .op(n11400) );
  nand2_1 U12142 ( .ip1(data_rd_mem[16]), .ip2(n12325), .op(n11399) );
  nand2_1 U12143 ( .ip1(n11400), .ip2(n11399), .op(n11570) );
  mux2_1 U12144 ( .ip1(\cache_data[0][16] ), .ip2(n11570), .s(n11415), .op(
        n6815) );
  nand2_1 U12145 ( .ip1(iCache_data_wr[17]), .ip2(n12323), .op(n11402) );
  nand2_1 U12146 ( .ip1(data_rd_mem[17]), .ip2(n12325), .op(n11401) );
  nand2_1 U12147 ( .ip1(n11402), .ip2(n11401), .op(n11571) );
  mux2_1 U12148 ( .ip1(\cache_data[0][17] ), .ip2(n11571), .s(n11415), .op(
        n6814) );
  nand2_1 U12149 ( .ip1(iCache_data_wr[18]), .ip2(n12323), .op(n11404) );
  nand2_1 U12150 ( .ip1(data_rd_mem[18]), .ip2(n12325), .op(n11403) );
  nand2_1 U12151 ( .ip1(n11404), .ip2(n11403), .op(n11572) );
  mux2_1 U12152 ( .ip1(\cache_data[0][18] ), .ip2(n11572), .s(n11415), .op(
        n6813) );
  nand2_1 U12153 ( .ip1(iCache_data_wr[19]), .ip2(n12323), .op(n11406) );
  nand2_1 U12154 ( .ip1(data_rd_mem[19]), .ip2(n12325), .op(n11405) );
  nand2_1 U12155 ( .ip1(n11406), .ip2(n11405), .op(n11573) );
  mux2_1 U12156 ( .ip1(\cache_data[0][19] ), .ip2(n11573), .s(n11415), .op(
        n6812) );
  nand2_1 U12157 ( .ip1(iCache_data_wr[20]), .ip2(n12323), .op(n11408) );
  nand2_1 U12158 ( .ip1(data_rd_mem[20]), .ip2(n12325), .op(n11407) );
  nand2_1 U12159 ( .ip1(n11408), .ip2(n11407), .op(n11574) );
  mux2_1 U12160 ( .ip1(\cache_data[0][20] ), .ip2(n11574), .s(n11415), .op(
        n6811) );
  nand2_1 U12161 ( .ip1(iCache_data_wr[21]), .ip2(n12323), .op(n11410) );
  nand2_1 U12162 ( .ip1(data_rd_mem[21]), .ip2(n12325), .op(n11409) );
  nand2_1 U12163 ( .ip1(n11410), .ip2(n11409), .op(n11575) );
  mux2_1 U12164 ( .ip1(\cache_data[0][21] ), .ip2(n11575), .s(n11415), .op(
        n6810) );
  nand2_1 U12165 ( .ip1(iCache_data_wr[22]), .ip2(n12323), .op(n11412) );
  nand2_1 U12166 ( .ip1(data_rd_mem[22]), .ip2(n12325), .op(n11411) );
  nand2_1 U12167 ( .ip1(n11412), .ip2(n11411), .op(n11576) );
  mux2_1 U12168 ( .ip1(\cache_data[0][22] ), .ip2(n11576), .s(n11415), .op(
        n6809) );
  nand2_1 U12169 ( .ip1(iCache_data_wr[23]), .ip2(n12323), .op(n11414) );
  nand2_1 U12170 ( .ip1(data_rd_mem[23]), .ip2(n12325), .op(n11413) );
  nand2_1 U12171 ( .ip1(n11414), .ip2(n11413), .op(n11577) );
  mux2_1 U12172 ( .ip1(\cache_data[0][23] ), .ip2(n11577), .s(n11415), .op(
        n6808) );
  nand2_1 U12173 ( .ip1(iCache_data_wr[24]), .ip2(n12323), .op(n11417) );
  nand2_1 U12174 ( .ip1(data_rd_mem[24]), .ip2(n12325), .op(n11416) );
  nand2_1 U12175 ( .ip1(n11417), .ip2(n11416), .op(n11578) );
  mux2_1 U12176 ( .ip1(\cache_data[0][24] ), .ip2(n11578), .s(n11432), .op(
        n6807) );
  nand2_1 U12177 ( .ip1(iCache_data_wr[25]), .ip2(n12323), .op(n11419) );
  nand2_1 U12178 ( .ip1(data_rd_mem[25]), .ip2(n12325), .op(n11418) );
  nand2_1 U12179 ( .ip1(n11419), .ip2(n11418), .op(n11580) );
  mux2_1 U12180 ( .ip1(\cache_data[0][25] ), .ip2(n11580), .s(n11432), .op(
        n6806) );
  nand2_1 U12181 ( .ip1(iCache_data_wr[26]), .ip2(n12323), .op(n11421) );
  nand2_1 U12182 ( .ip1(data_rd_mem[26]), .ip2(n12325), .op(n11420) );
  nand2_1 U12183 ( .ip1(n11421), .ip2(n11420), .op(n11581) );
  mux2_1 U12184 ( .ip1(\cache_data[0][26] ), .ip2(n11581), .s(n11432), .op(
        n6805) );
  nand2_1 U12185 ( .ip1(iCache_data_wr[27]), .ip2(n12323), .op(n11423) );
  nand2_1 U12186 ( .ip1(data_rd_mem[27]), .ip2(n12325), .op(n11422) );
  nand2_1 U12187 ( .ip1(n11423), .ip2(n11422), .op(n11582) );
  mux2_1 U12188 ( .ip1(\cache_data[0][27] ), .ip2(n11582), .s(n11432), .op(
        n6804) );
  nand2_1 U12189 ( .ip1(iCache_data_wr[28]), .ip2(n12323), .op(n11425) );
  nand2_1 U12190 ( .ip1(data_rd_mem[28]), .ip2(n12325), .op(n11424) );
  nand2_1 U12191 ( .ip1(n11425), .ip2(n11424), .op(n11583) );
  mux2_1 U12192 ( .ip1(\cache_data[0][28] ), .ip2(n11583), .s(n11432), .op(
        n6803) );
  nand2_1 U12193 ( .ip1(iCache_data_wr[29]), .ip2(n12323), .op(n11427) );
  nand2_1 U12194 ( .ip1(data_rd_mem[29]), .ip2(n12325), .op(n11426) );
  nand2_1 U12195 ( .ip1(n11427), .ip2(n11426), .op(n11584) );
  mux2_1 U12196 ( .ip1(\cache_data[0][29] ), .ip2(n11584), .s(n11432), .op(
        n6802) );
  nand2_1 U12197 ( .ip1(iCache_data_wr[30]), .ip2(n12323), .op(n11429) );
  nand2_1 U12198 ( .ip1(data_rd_mem[30]), .ip2(n12325), .op(n11428) );
  nand2_1 U12199 ( .ip1(n11429), .ip2(n11428), .op(n11585) );
  mux2_1 U12200 ( .ip1(\cache_data[0][30] ), .ip2(n11585), .s(n11432), .op(
        n6801) );
  nand2_1 U12201 ( .ip1(iCache_data_wr[31]), .ip2(n12323), .op(n11431) );
  nand2_1 U12202 ( .ip1(data_rd_mem[31]), .ip2(n12325), .op(n11430) );
  nand2_1 U12203 ( .ip1(n11431), .ip2(n11430), .op(n11587) );
  mux2_1 U12204 ( .ip1(\cache_data[0][31] ), .ip2(n11587), .s(n11432), .op(
        n6800) );
  nor3_1 U12205 ( .ip1(addr_resp[3]), .ip2(n11445), .ip3(n11446), .op(n11435)
         );
  nor3_1 U12206 ( .ip1(mem_data_cnt[3]), .ip2(n11433), .ip3(n11443), .op(
        n11434) );
  nor2_1 U12207 ( .ip1(n11435), .ip2(n11434), .op(n11606) );
  nor2_1 U12208 ( .ip1(n11606), .ip2(n8923), .op(n11436) );
  mux2_1 U12209 ( .ip1(\cache_data[0][32] ), .ip2(n11554), .s(n11436), .op(
        n6799) );
  mux2_1 U12210 ( .ip1(\cache_data[0][33] ), .ip2(n11555), .s(n11436), .op(
        n6798) );
  mux2_1 U12211 ( .ip1(\cache_data[0][34] ), .ip2(n11556), .s(n11436), .op(
        n6797) );
  mux2_1 U12212 ( .ip1(\cache_data[0][35] ), .ip2(n11557), .s(n11436), .op(
        n6796) );
  mux2_1 U12213 ( .ip1(\cache_data[0][36] ), .ip2(n11558), .s(n11436), .op(
        n6795) );
  mux2_1 U12214 ( .ip1(\cache_data[0][37] ), .ip2(n11559), .s(n11436), .op(
        n6794) );
  mux2_1 U12215 ( .ip1(\cache_data[0][38] ), .ip2(n11560), .s(n11436), .op(
        n6793) );
  mux2_1 U12216 ( .ip1(\cache_data[0][39] ), .ip2(n11561), .s(n11436), .op(
        n6792) );
  mux2_1 U12217 ( .ip1(\cache_data[0][40] ), .ip2(n11562), .s(n11436), .op(
        n6791) );
  buf_1 U12218 ( .ip(n11436), .op(n11437) );
  mux2_1 U12219 ( .ip1(\cache_data[0][41] ), .ip2(n11563), .s(n11437), .op(
        n6790) );
  mux2_1 U12220 ( .ip1(\cache_data[0][42] ), .ip2(n11564), .s(n11437), .op(
        n6789) );
  mux2_1 U12221 ( .ip1(\cache_data[0][43] ), .ip2(n11565), .s(n11436), .op(
        n6788) );
  mux2_1 U12222 ( .ip1(\cache_data[0][44] ), .ip2(n11566), .s(n11436), .op(
        n6787) );
  mux2_1 U12223 ( .ip1(\cache_data[0][45] ), .ip2(n11567), .s(n11437), .op(
        n6786) );
  mux2_1 U12224 ( .ip1(\cache_data[0][46] ), .ip2(n11568), .s(n11436), .op(
        n6785) );
  mux2_1 U12225 ( .ip1(\cache_data[0][47] ), .ip2(n11569), .s(n11436), .op(
        n6784) );
  mux2_1 U12226 ( .ip1(\cache_data[0][48] ), .ip2(n11570), .s(n11436), .op(
        n6783) );
  mux2_1 U12227 ( .ip1(\cache_data[0][49] ), .ip2(n11571), .s(n11436), .op(
        n6782) );
  mux2_1 U12228 ( .ip1(\cache_data[0][50] ), .ip2(n11572), .s(n11436), .op(
        n6781) );
  mux2_1 U12229 ( .ip1(\cache_data[0][51] ), .ip2(n11573), .s(n11436), .op(
        n6780) );
  mux2_1 U12230 ( .ip1(\cache_data[0][52] ), .ip2(n11574), .s(n11436), .op(
        n6779) );
  mux2_1 U12231 ( .ip1(\cache_data[0][53] ), .ip2(n11575), .s(n11436), .op(
        n6778) );
  mux2_1 U12232 ( .ip1(\cache_data[0][54] ), .ip2(n11576), .s(n11436), .op(
        n6777) );
  mux2_1 U12233 ( .ip1(\cache_data[0][55] ), .ip2(n11577), .s(n11436), .op(
        n6776) );
  mux2_1 U12234 ( .ip1(\cache_data[0][56] ), .ip2(n11578), .s(n11437), .op(
        n6775) );
  mux2_1 U12235 ( .ip1(\cache_data[0][57] ), .ip2(n11580), .s(n11437), .op(
        n6774) );
  mux2_1 U12236 ( .ip1(\cache_data[0][58] ), .ip2(n11581), .s(n11437), .op(
        n6773) );
  mux2_1 U12237 ( .ip1(\cache_data[0][59] ), .ip2(n11582), .s(n11437), .op(
        n6772) );
  mux2_1 U12238 ( .ip1(\cache_data[0][60] ), .ip2(n11583), .s(n11437), .op(
        n6771) );
  mux2_1 U12239 ( .ip1(\cache_data[0][61] ), .ip2(n11584), .s(n11437), .op(
        n6770) );
  mux2_1 U12240 ( .ip1(\cache_data[0][62] ), .ip2(n11585), .s(n11437), .op(
        n6769) );
  mux2_1 U12241 ( .ip1(\cache_data[0][63] ), .ip2(n11587), .s(n11437), .op(
        n6768) );
  nor3_1 U12242 ( .ip1(addr_resp[2]), .ip2(n11446), .ip3(n11444), .op(n11440)
         );
  nor3_1 U12243 ( .ip1(mem_data_cnt[2]), .ip2(n11438), .ip3(n11443), .op(
        n11439) );
  nor2_1 U12244 ( .ip1(n11440), .ip2(n11439), .op(n11609) );
  nor2_1 U12245 ( .ip1(n11609), .ip2(n8923), .op(n11441) );
  mux2_1 U12246 ( .ip1(\cache_data[0][64] ), .ip2(n11554), .s(n11441), .op(
        n6767) );
  mux2_1 U12247 ( .ip1(\cache_data[0][65] ), .ip2(n11555), .s(n11441), .op(
        n6766) );
  mux2_1 U12248 ( .ip1(\cache_data[0][66] ), .ip2(n11556), .s(n11441), .op(
        n6765) );
  mux2_1 U12249 ( .ip1(\cache_data[0][67] ), .ip2(n11557), .s(n11441), .op(
        n6764) );
  mux2_1 U12250 ( .ip1(\cache_data[0][68] ), .ip2(n11558), .s(n11441), .op(
        n6763) );
  mux2_1 U12251 ( .ip1(\cache_data[0][69] ), .ip2(n11559), .s(n11441), .op(
        n6762) );
  mux2_1 U12252 ( .ip1(\cache_data[0][70] ), .ip2(n11560), .s(n11441), .op(
        n6761) );
  mux2_1 U12253 ( .ip1(\cache_data[0][71] ), .ip2(n11561), .s(n11441), .op(
        n6760) );
  mux2_1 U12254 ( .ip1(\cache_data[0][72] ), .ip2(n11562), .s(n11441), .op(
        n6759) );
  buf_1 U12255 ( .ip(n11441), .op(n11442) );
  mux2_1 U12256 ( .ip1(\cache_data[0][73] ), .ip2(n11563), .s(n11442), .op(
        n6758) );
  mux2_1 U12257 ( .ip1(\cache_data[0][74] ), .ip2(n11564), .s(n11442), .op(
        n6757) );
  mux2_1 U12258 ( .ip1(\cache_data[0][75] ), .ip2(n11565), .s(n11441), .op(
        n6756) );
  mux2_1 U12259 ( .ip1(\cache_data[0][76] ), .ip2(n11566), .s(n11441), .op(
        n6755) );
  mux2_1 U12260 ( .ip1(\cache_data[0][77] ), .ip2(n11567), .s(n11442), .op(
        n6754) );
  mux2_1 U12261 ( .ip1(\cache_data[0][78] ), .ip2(n11568), .s(n11441), .op(
        n6753) );
  mux2_1 U12262 ( .ip1(\cache_data[0][79] ), .ip2(n11569), .s(n11441), .op(
        n6752) );
  mux2_1 U12263 ( .ip1(\cache_data[0][80] ), .ip2(n11570), .s(n11441), .op(
        n6751) );
  mux2_1 U12264 ( .ip1(\cache_data[0][81] ), .ip2(n11571), .s(n11441), .op(
        n6750) );
  mux2_1 U12265 ( .ip1(\cache_data[0][82] ), .ip2(n11572), .s(n11441), .op(
        n6749) );
  mux2_1 U12266 ( .ip1(\cache_data[0][83] ), .ip2(n11573), .s(n11441), .op(
        n6748) );
  mux2_1 U12267 ( .ip1(\cache_data[0][84] ), .ip2(n11574), .s(n11441), .op(
        n6747) );
  mux2_1 U12268 ( .ip1(\cache_data[0][85] ), .ip2(n11575), .s(n11441), .op(
        n6746) );
  mux2_1 U12269 ( .ip1(\cache_data[0][86] ), .ip2(n11576), .s(n11441), .op(
        n6745) );
  mux2_1 U12270 ( .ip1(\cache_data[0][87] ), .ip2(n11577), .s(n11441), .op(
        n6744) );
  mux2_1 U12271 ( .ip1(\cache_data[0][88] ), .ip2(n11578), .s(n11442), .op(
        n6743) );
  mux2_1 U12272 ( .ip1(\cache_data[0][89] ), .ip2(n11580), .s(n11442), .op(
        n6742) );
  mux2_1 U12273 ( .ip1(\cache_data[0][90] ), .ip2(n11581), .s(n11442), .op(
        n6741) );
  mux2_1 U12274 ( .ip1(\cache_data[0][91] ), .ip2(n11582), .s(n11442), .op(
        n6740) );
  mux2_1 U12275 ( .ip1(\cache_data[0][92] ), .ip2(n11583), .s(n11442), .op(
        n6739) );
  mux2_1 U12276 ( .ip1(\cache_data[0][93] ), .ip2(n11584), .s(n11442), .op(
        n6738) );
  mux2_1 U12277 ( .ip1(\cache_data[0][94] ), .ip2(n11585), .s(n11442), .op(
        n6737) );
  mux2_1 U12278 ( .ip1(\cache_data[0][95] ), .ip2(n11587), .s(n11442), .op(
        n6736) );
  inv_1 U12279 ( .ip(n11443), .op(n11447) );
  nor3_1 U12280 ( .ip1(n11446), .ip2(n11445), .ip3(n11444), .op(n11448) );
  or2_1 U12281 ( .ip1(n11447), .ip2(n11448), .op(n11450) );
  or2_1 U12282 ( .ip1(N3698), .ip2(n11448), .op(n11449) );
  nand2_1 U12283 ( .ip1(n11450), .ip2(n11449), .op(n11613) );
  nor2_1 U12284 ( .ip1(n11613), .ip2(n8923), .op(n11451) );
  mux2_1 U12285 ( .ip1(\cache_data[0][96] ), .ip2(n11554), .s(n11451), .op(
        n6735) );
  mux2_1 U12286 ( .ip1(\cache_data[0][97] ), .ip2(n11555), .s(n11451), .op(
        n6734) );
  mux2_1 U12287 ( .ip1(\cache_data[0][98] ), .ip2(n11556), .s(n11451), .op(
        n6733) );
  mux2_1 U12288 ( .ip1(\cache_data[0][99] ), .ip2(n11557), .s(n11451), .op(
        n6732) );
  mux2_1 U12289 ( .ip1(\cache_data[0][100] ), .ip2(n11558), .s(n11451), .op(
        n6731) );
  mux2_1 U12290 ( .ip1(\cache_data[0][101] ), .ip2(n11559), .s(n11451), .op(
        n6730) );
  mux2_1 U12291 ( .ip1(\cache_data[0][102] ), .ip2(n11560), .s(n11451), .op(
        n6729) );
  mux2_1 U12292 ( .ip1(\cache_data[0][103] ), .ip2(n11561), .s(n11451), .op(
        n6728) );
  mux2_1 U12293 ( .ip1(\cache_data[0][104] ), .ip2(n11562), .s(n11451), .op(
        n6727) );
  buf_1 U12294 ( .ip(n11451), .op(n11452) );
  mux2_1 U12295 ( .ip1(\cache_data[0][105] ), .ip2(n11563), .s(n11452), .op(
        n6726) );
  mux2_1 U12296 ( .ip1(\cache_data[0][106] ), .ip2(n11564), .s(n11452), .op(
        n6725) );
  mux2_1 U12297 ( .ip1(\cache_data[0][107] ), .ip2(n11565), .s(n11451), .op(
        n6724) );
  mux2_1 U12298 ( .ip1(\cache_data[0][108] ), .ip2(n11566), .s(n11451), .op(
        n6723) );
  mux2_1 U12299 ( .ip1(\cache_data[0][109] ), .ip2(n11567), .s(n11452), .op(
        n6722) );
  mux2_1 U12300 ( .ip1(\cache_data[0][110] ), .ip2(n11568), .s(n11451), .op(
        n6721) );
  mux2_1 U12301 ( .ip1(\cache_data[0][111] ), .ip2(n11569), .s(n11451), .op(
        n6720) );
  mux2_1 U12302 ( .ip1(\cache_data[0][112] ), .ip2(n11570), .s(n11451), .op(
        n6719) );
  mux2_1 U12303 ( .ip1(\cache_data[0][113] ), .ip2(n11571), .s(n11451), .op(
        n6718) );
  mux2_1 U12304 ( .ip1(\cache_data[0][114] ), .ip2(n11572), .s(n11451), .op(
        n6717) );
  mux2_1 U12305 ( .ip1(\cache_data[0][115] ), .ip2(n11573), .s(n11451), .op(
        n6716) );
  mux2_1 U12306 ( .ip1(\cache_data[0][116] ), .ip2(n11574), .s(n11451), .op(
        n6715) );
  mux2_1 U12307 ( .ip1(\cache_data[0][117] ), .ip2(n11575), .s(n11451), .op(
        n6714) );
  mux2_1 U12308 ( .ip1(\cache_data[0][118] ), .ip2(n11576), .s(n11451), .op(
        n6713) );
  mux2_1 U12309 ( .ip1(\cache_data[0][119] ), .ip2(n11577), .s(n11451), .op(
        n6712) );
  mux2_1 U12310 ( .ip1(\cache_data[0][120] ), .ip2(n11578), .s(n11452), .op(
        n6711) );
  mux2_1 U12311 ( .ip1(\cache_data[0][121] ), .ip2(n11580), .s(n11452), .op(
        n6710) );
  mux2_1 U12312 ( .ip1(\cache_data[0][122] ), .ip2(n11581), .s(n11452), .op(
        n6709) );
  mux2_1 U12313 ( .ip1(\cache_data[0][123] ), .ip2(n11582), .s(n11452), .op(
        n6708) );
  mux2_1 U12314 ( .ip1(\cache_data[0][124] ), .ip2(n11583), .s(n11452), .op(
        n6707) );
  mux2_1 U12315 ( .ip1(\cache_data[0][125] ), .ip2(n11584), .s(n11452), .op(
        n6706) );
  mux2_1 U12316 ( .ip1(\cache_data[0][126] ), .ip2(n11585), .s(n11452), .op(
        n6705) );
  mux2_1 U12317 ( .ip1(\cache_data[0][127] ), .ip2(n11587), .s(n11452), .op(
        n6704) );
  nor2_1 U12318 ( .ip1(n11603), .ip2(n11459), .op(n11453) );
  mux2_1 U12319 ( .ip1(\cache_data[1][0] ), .ip2(n11554), .s(n11453), .op(
        n6703) );
  mux2_1 U12320 ( .ip1(\cache_data[1][1] ), .ip2(n11555), .s(n11453), .op(
        n6702) );
  mux2_1 U12321 ( .ip1(\cache_data[1][2] ), .ip2(n11556), .s(n11453), .op(
        n6701) );
  mux2_1 U12322 ( .ip1(\cache_data[1][3] ), .ip2(n11557), .s(n11453), .op(
        n6700) );
  mux2_1 U12323 ( .ip1(\cache_data[1][4] ), .ip2(n11558), .s(n11453), .op(
        n6699) );
  mux2_1 U12324 ( .ip1(\cache_data[1][5] ), .ip2(n11559), .s(n11453), .op(
        n6698) );
  mux2_1 U12325 ( .ip1(\cache_data[1][6] ), .ip2(n11560), .s(n11453), .op(
        n6697) );
  mux2_1 U12326 ( .ip1(\cache_data[1][7] ), .ip2(n11561), .s(n11453), .op(
        n6696) );
  mux2_1 U12327 ( .ip1(\cache_data[1][8] ), .ip2(n11562), .s(n11453), .op(
        n6695) );
  buf_1 U12328 ( .ip(n11453), .op(n11454) );
  mux2_1 U12329 ( .ip1(\cache_data[1][9] ), .ip2(n11563), .s(n11454), .op(
        n6694) );
  mux2_1 U12330 ( .ip1(\cache_data[1][10] ), .ip2(n11564), .s(n11454), .op(
        n6693) );
  mux2_1 U12331 ( .ip1(\cache_data[1][11] ), .ip2(n11565), .s(n11453), .op(
        n6692) );
  mux2_1 U12332 ( .ip1(\cache_data[1][12] ), .ip2(n11566), .s(n11453), .op(
        n6691) );
  mux2_1 U12333 ( .ip1(\cache_data[1][13] ), .ip2(n11567), .s(n11454), .op(
        n6690) );
  mux2_1 U12334 ( .ip1(\cache_data[1][14] ), .ip2(n11568), .s(n11453), .op(
        n6689) );
  mux2_1 U12335 ( .ip1(\cache_data[1][15] ), .ip2(n11569), .s(n11453), .op(
        n6688) );
  mux2_1 U12336 ( .ip1(\cache_data[1][16] ), .ip2(n11570), .s(n11453), .op(
        n6687) );
  mux2_1 U12337 ( .ip1(\cache_data[1][17] ), .ip2(n11571), .s(n11453), .op(
        n6686) );
  mux2_1 U12338 ( .ip1(\cache_data[1][18] ), .ip2(n11572), .s(n11453), .op(
        n6685) );
  mux2_1 U12339 ( .ip1(\cache_data[1][19] ), .ip2(n11573), .s(n11453), .op(
        n6684) );
  mux2_1 U12340 ( .ip1(\cache_data[1][20] ), .ip2(n11574), .s(n11453), .op(
        n6683) );
  mux2_1 U12341 ( .ip1(\cache_data[1][21] ), .ip2(n11575), .s(n11453), .op(
        n6682) );
  mux2_1 U12342 ( .ip1(\cache_data[1][22] ), .ip2(n11576), .s(n11453), .op(
        n6681) );
  mux2_1 U12343 ( .ip1(\cache_data[1][23] ), .ip2(n11577), .s(n11453), .op(
        n6680) );
  mux2_1 U12344 ( .ip1(\cache_data[1][24] ), .ip2(n11578), .s(n11454), .op(
        n6679) );
  mux2_1 U12345 ( .ip1(\cache_data[1][25] ), .ip2(n11580), .s(n11454), .op(
        n6678) );
  mux2_1 U12346 ( .ip1(\cache_data[1][26] ), .ip2(n11581), .s(n11454), .op(
        n6677) );
  mux2_1 U12347 ( .ip1(\cache_data[1][27] ), .ip2(n11582), .s(n11454), .op(
        n6676) );
  mux2_1 U12348 ( .ip1(\cache_data[1][28] ), .ip2(n11583), .s(n11454), .op(
        n6675) );
  mux2_1 U12349 ( .ip1(\cache_data[1][29] ), .ip2(n11584), .s(n11454), .op(
        n6674) );
  mux2_1 U12350 ( .ip1(\cache_data[1][30] ), .ip2(n11585), .s(n11454), .op(
        n6673) );
  mux2_1 U12351 ( .ip1(\cache_data[1][31] ), .ip2(n11587), .s(n11454), .op(
        n6672) );
  nor2_1 U12352 ( .ip1(n11606), .ip2(n11459), .op(n11455) );
  mux2_1 U12353 ( .ip1(\cache_data[1][32] ), .ip2(n11554), .s(n11455), .op(
        n6671) );
  mux2_1 U12354 ( .ip1(\cache_data[1][33] ), .ip2(n11555), .s(n11455), .op(
        n6670) );
  mux2_1 U12355 ( .ip1(\cache_data[1][34] ), .ip2(n11556), .s(n11455), .op(
        n6669) );
  mux2_1 U12356 ( .ip1(\cache_data[1][35] ), .ip2(n11557), .s(n11455), .op(
        n6668) );
  mux2_1 U12357 ( .ip1(\cache_data[1][36] ), .ip2(n11558), .s(n11455), .op(
        n6667) );
  mux2_1 U12358 ( .ip1(\cache_data[1][37] ), .ip2(n11559), .s(n11455), .op(
        n6666) );
  mux2_1 U12359 ( .ip1(\cache_data[1][38] ), .ip2(n11560), .s(n11455), .op(
        n6665) );
  mux2_1 U12360 ( .ip1(\cache_data[1][39] ), .ip2(n11561), .s(n11455), .op(
        n6664) );
  mux2_1 U12361 ( .ip1(\cache_data[1][40] ), .ip2(n11562), .s(n11455), .op(
        n6663) );
  buf_1 U12362 ( .ip(n11455), .op(n11456) );
  mux2_1 U12363 ( .ip1(\cache_data[1][41] ), .ip2(n11563), .s(n11456), .op(
        n6662) );
  mux2_1 U12364 ( .ip1(\cache_data[1][42] ), .ip2(n11564), .s(n11456), .op(
        n6661) );
  mux2_1 U12365 ( .ip1(\cache_data[1][43] ), .ip2(n11565), .s(n11455), .op(
        n6660) );
  mux2_1 U12366 ( .ip1(\cache_data[1][44] ), .ip2(n11566), .s(n11455), .op(
        n6659) );
  mux2_1 U12367 ( .ip1(\cache_data[1][45] ), .ip2(n11567), .s(n11456), .op(
        n6658) );
  mux2_1 U12368 ( .ip1(\cache_data[1][46] ), .ip2(n11568), .s(n11455), .op(
        n6657) );
  mux2_1 U12369 ( .ip1(\cache_data[1][47] ), .ip2(n11569), .s(n11455), .op(
        n6656) );
  mux2_1 U12370 ( .ip1(\cache_data[1][48] ), .ip2(n11570), .s(n11455), .op(
        n6655) );
  mux2_1 U12371 ( .ip1(\cache_data[1][49] ), .ip2(n11571), .s(n11455), .op(
        n6654) );
  mux2_1 U12372 ( .ip1(\cache_data[1][50] ), .ip2(n11572), .s(n11455), .op(
        n6653) );
  mux2_1 U12373 ( .ip1(\cache_data[1][51] ), .ip2(n11573), .s(n11455), .op(
        n6652) );
  mux2_1 U12374 ( .ip1(\cache_data[1][52] ), .ip2(n11574), .s(n11455), .op(
        n6651) );
  mux2_1 U12375 ( .ip1(\cache_data[1][53] ), .ip2(n11575), .s(n11455), .op(
        n6650) );
  mux2_1 U12376 ( .ip1(\cache_data[1][54] ), .ip2(n11576), .s(n11455), .op(
        n6649) );
  mux2_1 U12377 ( .ip1(\cache_data[1][55] ), .ip2(n11577), .s(n11455), .op(
        n6648) );
  mux2_1 U12378 ( .ip1(\cache_data[1][56] ), .ip2(n11578), .s(n11456), .op(
        n6647) );
  mux2_1 U12379 ( .ip1(\cache_data[1][57] ), .ip2(n11580), .s(n11456), .op(
        n6646) );
  mux2_1 U12380 ( .ip1(\cache_data[1][58] ), .ip2(n11581), .s(n11456), .op(
        n6645) );
  mux2_1 U12381 ( .ip1(\cache_data[1][59] ), .ip2(n11582), .s(n11456), .op(
        n6644) );
  mux2_1 U12382 ( .ip1(\cache_data[1][60] ), .ip2(n11583), .s(n11456), .op(
        n6643) );
  mux2_1 U12383 ( .ip1(\cache_data[1][61] ), .ip2(n11584), .s(n11456), .op(
        n6642) );
  mux2_1 U12384 ( .ip1(\cache_data[1][62] ), .ip2(n11585), .s(n11456), .op(
        n6641) );
  mux2_1 U12385 ( .ip1(\cache_data[1][63] ), .ip2(n11587), .s(n11456), .op(
        n6640) );
  nor2_1 U12386 ( .ip1(n11609), .ip2(n11459), .op(n11457) );
  mux2_1 U12387 ( .ip1(\cache_data[1][64] ), .ip2(n11554), .s(n11457), .op(
        n6639) );
  mux2_1 U12388 ( .ip1(\cache_data[1][65] ), .ip2(n11555), .s(n11457), .op(
        n6638) );
  mux2_1 U12389 ( .ip1(\cache_data[1][66] ), .ip2(n11556), .s(n11457), .op(
        n6637) );
  mux2_1 U12390 ( .ip1(\cache_data[1][67] ), .ip2(n11557), .s(n11457), .op(
        n6636) );
  mux2_1 U12391 ( .ip1(\cache_data[1][68] ), .ip2(n11558), .s(n11457), .op(
        n6635) );
  mux2_1 U12392 ( .ip1(\cache_data[1][69] ), .ip2(n11559), .s(n11457), .op(
        n6634) );
  mux2_1 U12393 ( .ip1(\cache_data[1][70] ), .ip2(n11560), .s(n11457), .op(
        n6633) );
  mux2_1 U12394 ( .ip1(\cache_data[1][71] ), .ip2(n11561), .s(n11457), .op(
        n6632) );
  mux2_1 U12395 ( .ip1(\cache_data[1][72] ), .ip2(n11562), .s(n11457), .op(
        n6631) );
  buf_1 U12396 ( .ip(n11457), .op(n11458) );
  mux2_1 U12397 ( .ip1(\cache_data[1][73] ), .ip2(n11563), .s(n11458), .op(
        n6630) );
  mux2_1 U12398 ( .ip1(\cache_data[1][74] ), .ip2(n11564), .s(n11458), .op(
        n6629) );
  mux2_1 U12399 ( .ip1(\cache_data[1][75] ), .ip2(n11565), .s(n11457), .op(
        n6628) );
  mux2_1 U12400 ( .ip1(\cache_data[1][76] ), .ip2(n11566), .s(n11457), .op(
        n6627) );
  mux2_1 U12401 ( .ip1(\cache_data[1][77] ), .ip2(n11567), .s(n11458), .op(
        n6626) );
  mux2_1 U12402 ( .ip1(\cache_data[1][78] ), .ip2(n11568), .s(n11457), .op(
        n6625) );
  mux2_1 U12403 ( .ip1(\cache_data[1][79] ), .ip2(n11569), .s(n11457), .op(
        n6624) );
  mux2_1 U12404 ( .ip1(\cache_data[1][80] ), .ip2(n11570), .s(n11457), .op(
        n6623) );
  mux2_1 U12405 ( .ip1(\cache_data[1][81] ), .ip2(n11571), .s(n11457), .op(
        n6622) );
  mux2_1 U12406 ( .ip1(\cache_data[1][82] ), .ip2(n11572), .s(n11457), .op(
        n6621) );
  mux2_1 U12407 ( .ip1(\cache_data[1][83] ), .ip2(n11573), .s(n11457), .op(
        n6620) );
  mux2_1 U12408 ( .ip1(\cache_data[1][84] ), .ip2(n11574), .s(n11457), .op(
        n6619) );
  mux2_1 U12409 ( .ip1(\cache_data[1][85] ), .ip2(n11575), .s(n11457), .op(
        n6618) );
  mux2_1 U12410 ( .ip1(\cache_data[1][86] ), .ip2(n11576), .s(n11457), .op(
        n6617) );
  mux2_1 U12411 ( .ip1(\cache_data[1][87] ), .ip2(n11577), .s(n11457), .op(
        n6616) );
  mux2_1 U12412 ( .ip1(\cache_data[1][88] ), .ip2(n11578), .s(n11458), .op(
        n6615) );
  mux2_1 U12413 ( .ip1(\cache_data[1][89] ), .ip2(n11580), .s(n11458), .op(
        n6614) );
  mux2_1 U12414 ( .ip1(\cache_data[1][90] ), .ip2(n11581), .s(n11458), .op(
        n6613) );
  mux2_1 U12415 ( .ip1(\cache_data[1][91] ), .ip2(n11582), .s(n11458), .op(
        n6612) );
  mux2_1 U12416 ( .ip1(\cache_data[1][92] ), .ip2(n11583), .s(n11458), .op(
        n6611) );
  mux2_1 U12417 ( .ip1(\cache_data[1][93] ), .ip2(n11584), .s(n11458), .op(
        n6610) );
  mux2_1 U12418 ( .ip1(\cache_data[1][94] ), .ip2(n11585), .s(n11458), .op(
        n6609) );
  mux2_1 U12419 ( .ip1(\cache_data[1][95] ), .ip2(n11587), .s(n11458), .op(
        n6608) );
  nor2_1 U12420 ( .ip1(n11613), .ip2(n11459), .op(n11460) );
  mux2_1 U12421 ( .ip1(\cache_data[1][96] ), .ip2(n11554), .s(n11460), .op(
        n6607) );
  mux2_1 U12422 ( .ip1(\cache_data[1][97] ), .ip2(n11555), .s(n11460), .op(
        n6606) );
  mux2_1 U12423 ( .ip1(\cache_data[1][98] ), .ip2(n11556), .s(n11460), .op(
        n6605) );
  mux2_1 U12424 ( .ip1(\cache_data[1][99] ), .ip2(n11557), .s(n11460), .op(
        n6604) );
  mux2_1 U12425 ( .ip1(\cache_data[1][100] ), .ip2(n11558), .s(n11460), .op(
        n6603) );
  mux2_1 U12426 ( .ip1(\cache_data[1][101] ), .ip2(n11559), .s(n11460), .op(
        n6602) );
  mux2_1 U12427 ( .ip1(\cache_data[1][102] ), .ip2(n11560), .s(n11460), .op(
        n6601) );
  mux2_1 U12428 ( .ip1(\cache_data[1][103] ), .ip2(n11561), .s(n11460), .op(
        n6600) );
  mux2_1 U12429 ( .ip1(\cache_data[1][104] ), .ip2(n11562), .s(n11460), .op(
        n6599) );
  buf_1 U12430 ( .ip(n11460), .op(n11461) );
  mux2_1 U12431 ( .ip1(\cache_data[1][105] ), .ip2(n11563), .s(n11461), .op(
        n6598) );
  mux2_1 U12432 ( .ip1(\cache_data[1][106] ), .ip2(n11564), .s(n11461), .op(
        n6597) );
  mux2_1 U12433 ( .ip1(\cache_data[1][107] ), .ip2(n11565), .s(n11460), .op(
        n6596) );
  mux2_1 U12434 ( .ip1(\cache_data[1][108] ), .ip2(n11566), .s(n11460), .op(
        n6595) );
  mux2_1 U12435 ( .ip1(\cache_data[1][109] ), .ip2(n11567), .s(n11461), .op(
        n6594) );
  mux2_1 U12436 ( .ip1(\cache_data[1][110] ), .ip2(n11568), .s(n11460), .op(
        n6593) );
  mux2_1 U12437 ( .ip1(\cache_data[1][111] ), .ip2(n11569), .s(n11460), .op(
        n6592) );
  mux2_1 U12438 ( .ip1(\cache_data[1][112] ), .ip2(n11570), .s(n11460), .op(
        n6591) );
  mux2_1 U12439 ( .ip1(\cache_data[1][113] ), .ip2(n11571), .s(n11460), .op(
        n6590) );
  mux2_1 U12440 ( .ip1(\cache_data[1][114] ), .ip2(n11572), .s(n11460), .op(
        n6589) );
  mux2_1 U12441 ( .ip1(\cache_data[1][115] ), .ip2(n11573), .s(n11460), .op(
        n6588) );
  mux2_1 U12442 ( .ip1(\cache_data[1][116] ), .ip2(n11574), .s(n11460), .op(
        n6587) );
  mux2_1 U12443 ( .ip1(\cache_data[1][117] ), .ip2(n11575), .s(n11460), .op(
        n6586) );
  mux2_1 U12444 ( .ip1(\cache_data[1][118] ), .ip2(n11576), .s(n11460), .op(
        n6585) );
  mux2_1 U12445 ( .ip1(\cache_data[1][119] ), .ip2(n11577), .s(n11460), .op(
        n6584) );
  mux2_1 U12446 ( .ip1(\cache_data[1][120] ), .ip2(n11578), .s(n11461), .op(
        n6583) );
  mux2_1 U12447 ( .ip1(\cache_data[1][121] ), .ip2(n11580), .s(n11461), .op(
        n6582) );
  mux2_1 U12448 ( .ip1(\cache_data[1][122] ), .ip2(n11581), .s(n11461), .op(
        n6581) );
  mux2_1 U12449 ( .ip1(\cache_data[1][123] ), .ip2(n11582), .s(n11461), .op(
        n6580) );
  mux2_1 U12450 ( .ip1(\cache_data[1][124] ), .ip2(n11583), .s(n11461), .op(
        n6579) );
  mux2_1 U12451 ( .ip1(\cache_data[1][125] ), .ip2(n11584), .s(n11461), .op(
        n6578) );
  mux2_1 U12452 ( .ip1(\cache_data[1][126] ), .ip2(n11585), .s(n11461), .op(
        n6577) );
  mux2_1 U12453 ( .ip1(\cache_data[1][127] ), .ip2(n11587), .s(n11461), .op(
        n6576) );
  nor2_1 U12454 ( .ip1(n11603), .ip2(n8928), .op(n11462) );
  mux2_1 U12455 ( .ip1(\cache_data[2][0] ), .ip2(n11554), .s(n11462), .op(
        n6575) );
  mux2_1 U12456 ( .ip1(\cache_data[2][1] ), .ip2(n11555), .s(n11462), .op(
        n6574) );
  mux2_1 U12457 ( .ip1(\cache_data[2][2] ), .ip2(n11556), .s(n11462), .op(
        n6573) );
  mux2_1 U12458 ( .ip1(\cache_data[2][3] ), .ip2(n11557), .s(n11462), .op(
        n6572) );
  mux2_1 U12459 ( .ip1(\cache_data[2][4] ), .ip2(n11558), .s(n11462), .op(
        n6571) );
  mux2_1 U12460 ( .ip1(\cache_data[2][5] ), .ip2(n11559), .s(n11462), .op(
        n6570) );
  mux2_1 U12461 ( .ip1(\cache_data[2][6] ), .ip2(n11560), .s(n11462), .op(
        n6569) );
  mux2_1 U12462 ( .ip1(\cache_data[2][7] ), .ip2(n11561), .s(n11462), .op(
        n6568) );
  mux2_1 U12463 ( .ip1(\cache_data[2][8] ), .ip2(n11562), .s(n11462), .op(
        n6567) );
  buf_1 U12464 ( .ip(n11462), .op(n11463) );
  mux2_1 U12465 ( .ip1(\cache_data[2][9] ), .ip2(n11563), .s(n11463), .op(
        n6566) );
  mux2_1 U12466 ( .ip1(\cache_data[2][10] ), .ip2(n11564), .s(n11463), .op(
        n6565) );
  mux2_1 U12467 ( .ip1(\cache_data[2][11] ), .ip2(n11565), .s(n11462), .op(
        n6564) );
  mux2_1 U12468 ( .ip1(\cache_data[2][12] ), .ip2(n11566), .s(n11462), .op(
        n6563) );
  mux2_1 U12469 ( .ip1(\cache_data[2][13] ), .ip2(n11567), .s(n11463), .op(
        n6562) );
  mux2_1 U12470 ( .ip1(\cache_data[2][14] ), .ip2(n11568), .s(n11462), .op(
        n6561) );
  mux2_1 U12471 ( .ip1(\cache_data[2][15] ), .ip2(n11569), .s(n11462), .op(
        n6560) );
  mux2_1 U12472 ( .ip1(\cache_data[2][16] ), .ip2(n11570), .s(n11462), .op(
        n6559) );
  mux2_1 U12473 ( .ip1(\cache_data[2][17] ), .ip2(n11571), .s(n11462), .op(
        n6558) );
  mux2_1 U12474 ( .ip1(\cache_data[2][18] ), .ip2(n11572), .s(n11462), .op(
        n6557) );
  mux2_1 U12475 ( .ip1(\cache_data[2][19] ), .ip2(n11573), .s(n11462), .op(
        n6556) );
  mux2_1 U12476 ( .ip1(\cache_data[2][20] ), .ip2(n11574), .s(n11462), .op(
        n6555) );
  mux2_1 U12477 ( .ip1(\cache_data[2][21] ), .ip2(n11575), .s(n11462), .op(
        n6554) );
  mux2_1 U12478 ( .ip1(\cache_data[2][22] ), .ip2(n11576), .s(n11462), .op(
        n6553) );
  mux2_1 U12479 ( .ip1(\cache_data[2][23] ), .ip2(n11577), .s(n11462), .op(
        n6552) );
  mux2_1 U12480 ( .ip1(\cache_data[2][24] ), .ip2(n11578), .s(n11463), .op(
        n6551) );
  mux2_1 U12481 ( .ip1(\cache_data[2][25] ), .ip2(n11580), .s(n11463), .op(
        n6550) );
  mux2_1 U12482 ( .ip1(\cache_data[2][26] ), .ip2(n11581), .s(n11463), .op(
        n6549) );
  mux2_1 U12483 ( .ip1(\cache_data[2][27] ), .ip2(n11582), .s(n11463), .op(
        n6548) );
  mux2_1 U12484 ( .ip1(\cache_data[2][28] ), .ip2(n11583), .s(n11463), .op(
        n6547) );
  mux2_1 U12485 ( .ip1(\cache_data[2][29] ), .ip2(n11584), .s(n11463), .op(
        n6546) );
  mux2_1 U12486 ( .ip1(\cache_data[2][30] ), .ip2(n11585), .s(n11463), .op(
        n6545) );
  mux2_1 U12487 ( .ip1(\cache_data[2][31] ), .ip2(n11587), .s(n11463), .op(
        n6544) );
  nor2_1 U12488 ( .ip1(n11606), .ip2(n8928), .op(n11464) );
  mux2_1 U12489 ( .ip1(\cache_data[2][32] ), .ip2(n11554), .s(n11464), .op(
        n6543) );
  mux2_1 U12490 ( .ip1(\cache_data[2][33] ), .ip2(n11555), .s(n11464), .op(
        n6542) );
  mux2_1 U12491 ( .ip1(\cache_data[2][34] ), .ip2(n11556), .s(n11464), .op(
        n6541) );
  mux2_1 U12492 ( .ip1(\cache_data[2][35] ), .ip2(n11557), .s(n11464), .op(
        n6540) );
  mux2_1 U12493 ( .ip1(\cache_data[2][36] ), .ip2(n11558), .s(n11464), .op(
        n6539) );
  mux2_1 U12494 ( .ip1(\cache_data[2][37] ), .ip2(n11559), .s(n11464), .op(
        n6538) );
  mux2_1 U12495 ( .ip1(\cache_data[2][38] ), .ip2(n11560), .s(n11464), .op(
        n6537) );
  mux2_1 U12496 ( .ip1(\cache_data[2][39] ), .ip2(n11561), .s(n11464), .op(
        n6536) );
  mux2_1 U12497 ( .ip1(\cache_data[2][40] ), .ip2(n11562), .s(n11464), .op(
        n6535) );
  buf_1 U12498 ( .ip(n11464), .op(n11465) );
  mux2_1 U12499 ( .ip1(\cache_data[2][41] ), .ip2(n11563), .s(n11465), .op(
        n6534) );
  mux2_1 U12500 ( .ip1(\cache_data[2][42] ), .ip2(n11564), .s(n11465), .op(
        n6533) );
  mux2_1 U12501 ( .ip1(\cache_data[2][43] ), .ip2(n11565), .s(n11464), .op(
        n6532) );
  mux2_1 U12502 ( .ip1(\cache_data[2][44] ), .ip2(n11566), .s(n11464), .op(
        n6531) );
  mux2_1 U12503 ( .ip1(\cache_data[2][45] ), .ip2(n11567), .s(n11465), .op(
        n6530) );
  mux2_1 U12504 ( .ip1(\cache_data[2][46] ), .ip2(n11568), .s(n11464), .op(
        n6529) );
  mux2_1 U12505 ( .ip1(\cache_data[2][47] ), .ip2(n11569), .s(n11464), .op(
        n6528) );
  mux2_1 U12506 ( .ip1(\cache_data[2][48] ), .ip2(n11570), .s(n11464), .op(
        n6527) );
  mux2_1 U12507 ( .ip1(\cache_data[2][49] ), .ip2(n11571), .s(n11464), .op(
        n6526) );
  mux2_1 U12508 ( .ip1(\cache_data[2][50] ), .ip2(n11572), .s(n11464), .op(
        n6525) );
  mux2_1 U12509 ( .ip1(\cache_data[2][51] ), .ip2(n11573), .s(n11464), .op(
        n6524) );
  mux2_1 U12510 ( .ip1(\cache_data[2][52] ), .ip2(n11574), .s(n11464), .op(
        n6523) );
  mux2_1 U12511 ( .ip1(\cache_data[2][53] ), .ip2(n11575), .s(n11464), .op(
        n6522) );
  mux2_1 U12512 ( .ip1(\cache_data[2][54] ), .ip2(n11576), .s(n11464), .op(
        n6521) );
  mux2_1 U12513 ( .ip1(\cache_data[2][55] ), .ip2(n11577), .s(n11464), .op(
        n6520) );
  mux2_1 U12514 ( .ip1(\cache_data[2][56] ), .ip2(n11578), .s(n11465), .op(
        n6519) );
  mux2_1 U12515 ( .ip1(\cache_data[2][57] ), .ip2(n11580), .s(n11465), .op(
        n6518) );
  mux2_1 U12516 ( .ip1(\cache_data[2][58] ), .ip2(n11581), .s(n11465), .op(
        n6517) );
  mux2_1 U12517 ( .ip1(\cache_data[2][59] ), .ip2(n11582), .s(n11465), .op(
        n6516) );
  mux2_1 U12518 ( .ip1(\cache_data[2][60] ), .ip2(n11583), .s(n11465), .op(
        n6515) );
  mux2_1 U12519 ( .ip1(\cache_data[2][61] ), .ip2(n11584), .s(n11465), .op(
        n6514) );
  mux2_1 U12520 ( .ip1(\cache_data[2][62] ), .ip2(n11585), .s(n11465), .op(
        n6513) );
  mux2_1 U12521 ( .ip1(\cache_data[2][63] ), .ip2(n11587), .s(n11465), .op(
        n6512) );
  nor2_1 U12522 ( .ip1(n11609), .ip2(n8928), .op(n11466) );
  mux2_1 U12523 ( .ip1(\cache_data[2][64] ), .ip2(n11554), .s(n11466), .op(
        n6511) );
  mux2_1 U12524 ( .ip1(\cache_data[2][65] ), .ip2(n11555), .s(n11466), .op(
        n6510) );
  mux2_1 U12525 ( .ip1(\cache_data[2][66] ), .ip2(n11556), .s(n11466), .op(
        n6509) );
  mux2_1 U12526 ( .ip1(\cache_data[2][67] ), .ip2(n11557), .s(n11466), .op(
        n6508) );
  mux2_1 U12527 ( .ip1(\cache_data[2][68] ), .ip2(n11558), .s(n11466), .op(
        n6507) );
  mux2_1 U12528 ( .ip1(\cache_data[2][69] ), .ip2(n11559), .s(n11466), .op(
        n6506) );
  mux2_1 U12529 ( .ip1(\cache_data[2][70] ), .ip2(n11560), .s(n11466), .op(
        n6505) );
  mux2_1 U12530 ( .ip1(\cache_data[2][71] ), .ip2(n11561), .s(n11466), .op(
        n6504) );
  mux2_1 U12531 ( .ip1(\cache_data[2][72] ), .ip2(n11562), .s(n11466), .op(
        n6503) );
  buf_1 U12532 ( .ip(n11466), .op(n11467) );
  mux2_1 U12533 ( .ip1(\cache_data[2][73] ), .ip2(n11563), .s(n11467), .op(
        n6502) );
  mux2_1 U12534 ( .ip1(\cache_data[2][74] ), .ip2(n11564), .s(n11467), .op(
        n6501) );
  mux2_1 U12535 ( .ip1(\cache_data[2][75] ), .ip2(n11565), .s(n11466), .op(
        n6500) );
  mux2_1 U12536 ( .ip1(\cache_data[2][76] ), .ip2(n11566), .s(n11466), .op(
        n6499) );
  mux2_1 U12537 ( .ip1(\cache_data[2][77] ), .ip2(n11567), .s(n11467), .op(
        n6498) );
  mux2_1 U12538 ( .ip1(\cache_data[2][78] ), .ip2(n11568), .s(n11466), .op(
        n6497) );
  mux2_1 U12539 ( .ip1(\cache_data[2][79] ), .ip2(n11569), .s(n11466), .op(
        n6496) );
  mux2_1 U12540 ( .ip1(\cache_data[2][80] ), .ip2(n11570), .s(n11466), .op(
        n6495) );
  mux2_1 U12541 ( .ip1(\cache_data[2][81] ), .ip2(n11571), .s(n11466), .op(
        n6494) );
  mux2_1 U12542 ( .ip1(\cache_data[2][82] ), .ip2(n11572), .s(n11466), .op(
        n6493) );
  mux2_1 U12543 ( .ip1(\cache_data[2][83] ), .ip2(n11573), .s(n11466), .op(
        n6492) );
  mux2_1 U12544 ( .ip1(\cache_data[2][84] ), .ip2(n11574), .s(n11466), .op(
        n6491) );
  mux2_1 U12545 ( .ip1(\cache_data[2][85] ), .ip2(n11575), .s(n11466), .op(
        n6490) );
  mux2_1 U12546 ( .ip1(\cache_data[2][86] ), .ip2(n11576), .s(n11466), .op(
        n6489) );
  mux2_1 U12547 ( .ip1(\cache_data[2][87] ), .ip2(n11577), .s(n11466), .op(
        n6488) );
  mux2_1 U12548 ( .ip1(\cache_data[2][88] ), .ip2(n11578), .s(n11467), .op(
        n6487) );
  mux2_1 U12549 ( .ip1(\cache_data[2][89] ), .ip2(n11580), .s(n11467), .op(
        n6486) );
  mux2_1 U12550 ( .ip1(\cache_data[2][90] ), .ip2(n11581), .s(n11467), .op(
        n6485) );
  mux2_1 U12551 ( .ip1(\cache_data[2][91] ), .ip2(n11582), .s(n11467), .op(
        n6484) );
  mux2_1 U12552 ( .ip1(\cache_data[2][92] ), .ip2(n11583), .s(n11467), .op(
        n6483) );
  mux2_1 U12553 ( .ip1(\cache_data[2][93] ), .ip2(n11584), .s(n11467), .op(
        n6482) );
  mux2_1 U12554 ( .ip1(\cache_data[2][94] ), .ip2(n11585), .s(n11467), .op(
        n6481) );
  mux2_1 U12555 ( .ip1(\cache_data[2][95] ), .ip2(n11587), .s(n11467), .op(
        n6480) );
  nor2_1 U12556 ( .ip1(n11613), .ip2(n8928), .op(n11468) );
  mux2_1 U12557 ( .ip1(\cache_data[2][96] ), .ip2(n11554), .s(n11468), .op(
        n6479) );
  mux2_1 U12558 ( .ip1(\cache_data[2][97] ), .ip2(n11555), .s(n11468), .op(
        n6478) );
  mux2_1 U12559 ( .ip1(\cache_data[2][98] ), .ip2(n11556), .s(n11468), .op(
        n6477) );
  mux2_1 U12560 ( .ip1(\cache_data[2][99] ), .ip2(n11557), .s(n11468), .op(
        n6476) );
  mux2_1 U12561 ( .ip1(\cache_data[2][100] ), .ip2(n11558), .s(n11468), .op(
        n6475) );
  mux2_1 U12562 ( .ip1(\cache_data[2][101] ), .ip2(n11559), .s(n11468), .op(
        n6474) );
  mux2_1 U12563 ( .ip1(\cache_data[2][102] ), .ip2(n11560), .s(n11468), .op(
        n6473) );
  mux2_1 U12564 ( .ip1(\cache_data[2][103] ), .ip2(n11561), .s(n11468), .op(
        n6472) );
  mux2_1 U12565 ( .ip1(\cache_data[2][104] ), .ip2(n11562), .s(n11468), .op(
        n6471) );
  buf_1 U12566 ( .ip(n11468), .op(n11469) );
  mux2_1 U12567 ( .ip1(\cache_data[2][105] ), .ip2(n11563), .s(n11469), .op(
        n6470) );
  mux2_1 U12568 ( .ip1(\cache_data[2][106] ), .ip2(n11564), .s(n11469), .op(
        n6469) );
  mux2_1 U12569 ( .ip1(\cache_data[2][107] ), .ip2(n11565), .s(n11468), .op(
        n6468) );
  mux2_1 U12570 ( .ip1(\cache_data[2][108] ), .ip2(n11566), .s(n11468), .op(
        n6467) );
  mux2_1 U12571 ( .ip1(\cache_data[2][109] ), .ip2(n11567), .s(n11469), .op(
        n6466) );
  mux2_1 U12572 ( .ip1(\cache_data[2][110] ), .ip2(n11568), .s(n11468), .op(
        n6465) );
  mux2_1 U12573 ( .ip1(\cache_data[2][111] ), .ip2(n11569), .s(n11468), .op(
        n6464) );
  mux2_1 U12574 ( .ip1(\cache_data[2][112] ), .ip2(n11570), .s(n11468), .op(
        n6463) );
  mux2_1 U12575 ( .ip1(\cache_data[2][113] ), .ip2(n11571), .s(n11468), .op(
        n6462) );
  mux2_1 U12576 ( .ip1(\cache_data[2][114] ), .ip2(n11572), .s(n11468), .op(
        n6461) );
  mux2_1 U12577 ( .ip1(\cache_data[2][115] ), .ip2(n11573), .s(n11468), .op(
        n6460) );
  mux2_1 U12578 ( .ip1(\cache_data[2][116] ), .ip2(n11574), .s(n11468), .op(
        n6459) );
  mux2_1 U12579 ( .ip1(\cache_data[2][117] ), .ip2(n11575), .s(n11468), .op(
        n6458) );
  mux2_1 U12580 ( .ip1(\cache_data[2][118] ), .ip2(n11576), .s(n11468), .op(
        n6457) );
  mux2_1 U12581 ( .ip1(\cache_data[2][119] ), .ip2(n11577), .s(n11468), .op(
        n6456) );
  mux2_1 U12582 ( .ip1(\cache_data[2][120] ), .ip2(n11578), .s(n11469), .op(
        n6455) );
  mux2_1 U12583 ( .ip1(\cache_data[2][121] ), .ip2(n11580), .s(n11469), .op(
        n6454) );
  mux2_1 U12584 ( .ip1(\cache_data[2][122] ), .ip2(n11581), .s(n11469), .op(
        n6453) );
  mux2_1 U12585 ( .ip1(\cache_data[2][123] ), .ip2(n11582), .s(n11469), .op(
        n6452) );
  mux2_1 U12586 ( .ip1(\cache_data[2][124] ), .ip2(n11583), .s(n11469), .op(
        n6451) );
  mux2_1 U12587 ( .ip1(\cache_data[2][125] ), .ip2(n11584), .s(n11469), .op(
        n6450) );
  mux2_1 U12588 ( .ip1(\cache_data[2][126] ), .ip2(n11585), .s(n11469), .op(
        n6449) );
  mux2_1 U12589 ( .ip1(\cache_data[2][127] ), .ip2(n11587), .s(n11469), .op(
        n6448) );
  nor2_1 U12590 ( .ip1(n11603), .ip2(n11476), .op(n11470) );
  mux2_1 U12591 ( .ip1(\cache_data[3][0] ), .ip2(n11554), .s(n11470), .op(
        n6447) );
  mux2_1 U12592 ( .ip1(\cache_data[3][1] ), .ip2(n11555), .s(n11470), .op(
        n6446) );
  mux2_1 U12593 ( .ip1(\cache_data[3][2] ), .ip2(n11556), .s(n11470), .op(
        n6445) );
  mux2_1 U12594 ( .ip1(\cache_data[3][3] ), .ip2(n11557), .s(n11470), .op(
        n6444) );
  mux2_1 U12595 ( .ip1(\cache_data[3][4] ), .ip2(n11558), .s(n11470), .op(
        n6443) );
  mux2_1 U12596 ( .ip1(\cache_data[3][5] ), .ip2(n11559), .s(n11470), .op(
        n6442) );
  mux2_1 U12597 ( .ip1(\cache_data[3][6] ), .ip2(n11560), .s(n11470), .op(
        n6441) );
  mux2_1 U12598 ( .ip1(\cache_data[3][7] ), .ip2(n11561), .s(n11470), .op(
        n6440) );
  mux2_1 U12599 ( .ip1(\cache_data[3][8] ), .ip2(n11562), .s(n11470), .op(
        n6439) );
  mux2_1 U12600 ( .ip1(\cache_data[3][9] ), .ip2(n11563), .s(n11470), .op(
        n6438) );
  mux2_1 U12601 ( .ip1(\cache_data[3][10] ), .ip2(n11564), .s(n11470), .op(
        n6437) );
  mux2_1 U12602 ( .ip1(\cache_data[3][11] ), .ip2(n11565), .s(n11470), .op(
        n6436) );
  mux2_1 U12603 ( .ip1(\cache_data[3][12] ), .ip2(n11566), .s(n11470), .op(
        n6435) );
  mux2_1 U12604 ( .ip1(\cache_data[3][13] ), .ip2(n11567), .s(n11470), .op(
        n6434) );
  mux2_1 U12605 ( .ip1(\cache_data[3][14] ), .ip2(n11568), .s(n11470), .op(
        n6433) );
  mux2_1 U12606 ( .ip1(\cache_data[3][15] ), .ip2(n11569), .s(n11470), .op(
        n6432) );
  mux2_1 U12607 ( .ip1(\cache_data[3][16] ), .ip2(n11570), .s(n11470), .op(
        n6431) );
  mux2_1 U12608 ( .ip1(\cache_data[3][17] ), .ip2(n11571), .s(n11470), .op(
        n6430) );
  mux2_1 U12609 ( .ip1(\cache_data[3][18] ), .ip2(n11572), .s(n11470), .op(
        n6429) );
  buf_1 U12610 ( .ip(n11470), .op(n11471) );
  mux2_1 U12611 ( .ip1(\cache_data[3][19] ), .ip2(n11573), .s(n11471), .op(
        n6428) );
  mux2_1 U12612 ( .ip1(\cache_data[3][20] ), .ip2(n11574), .s(n11471), .op(
        n6427) );
  mux2_1 U12613 ( .ip1(\cache_data[3][21] ), .ip2(n11575), .s(n11471), .op(
        n6426) );
  mux2_1 U12614 ( .ip1(\cache_data[3][22] ), .ip2(n11576), .s(n11471), .op(
        n6425) );
  mux2_1 U12615 ( .ip1(\cache_data[3][23] ), .ip2(n11577), .s(n11471), .op(
        n6424) );
  mux2_1 U12616 ( .ip1(\cache_data[3][24] ), .ip2(n11578), .s(n11470), .op(
        n6423) );
  mux2_1 U12617 ( .ip1(\cache_data[3][25] ), .ip2(n11580), .s(n11470), .op(
        n6422) );
  mux2_1 U12618 ( .ip1(\cache_data[3][26] ), .ip2(n11581), .s(n11471), .op(
        n6421) );
  mux2_1 U12619 ( .ip1(\cache_data[3][27] ), .ip2(n11582), .s(n11471), .op(
        n6420) );
  mux2_1 U12620 ( .ip1(\cache_data[3][28] ), .ip2(n11583), .s(n11471), .op(
        n6419) );
  mux2_1 U12621 ( .ip1(\cache_data[3][29] ), .ip2(n11584), .s(n11471), .op(
        n6418) );
  mux2_1 U12622 ( .ip1(\cache_data[3][30] ), .ip2(n11585), .s(n11471), .op(
        n6417) );
  mux2_1 U12623 ( .ip1(\cache_data[3][31] ), .ip2(n11587), .s(n11471), .op(
        n6416) );
  nor2_1 U12624 ( .ip1(n11606), .ip2(n11476), .op(n11472) );
  mux2_1 U12625 ( .ip1(\cache_data[3][32] ), .ip2(n11554), .s(n11472), .op(
        n6415) );
  mux2_1 U12626 ( .ip1(\cache_data[3][33] ), .ip2(n11555), .s(n11472), .op(
        n6414) );
  mux2_1 U12627 ( .ip1(\cache_data[3][34] ), .ip2(n11556), .s(n11472), .op(
        n6413) );
  mux2_1 U12628 ( .ip1(\cache_data[3][35] ), .ip2(n11557), .s(n11472), .op(
        n6412) );
  mux2_1 U12629 ( .ip1(\cache_data[3][36] ), .ip2(n11558), .s(n11472), .op(
        n6411) );
  mux2_1 U12630 ( .ip1(\cache_data[3][37] ), .ip2(n11559), .s(n11472), .op(
        n6410) );
  mux2_1 U12631 ( .ip1(\cache_data[3][38] ), .ip2(n11560), .s(n11472), .op(
        n6409) );
  mux2_1 U12632 ( .ip1(\cache_data[3][39] ), .ip2(n11561), .s(n11472), .op(
        n6408) );
  mux2_1 U12633 ( .ip1(\cache_data[3][40] ), .ip2(n11562), .s(n11472), .op(
        n6407) );
  mux2_1 U12634 ( .ip1(\cache_data[3][41] ), .ip2(n11563), .s(n11472), .op(
        n6406) );
  mux2_1 U12635 ( .ip1(\cache_data[3][42] ), .ip2(n11564), .s(n11472), .op(
        n6405) );
  mux2_1 U12636 ( .ip1(\cache_data[3][43] ), .ip2(n11565), .s(n11472), .op(
        n6404) );
  mux2_1 U12637 ( .ip1(\cache_data[3][44] ), .ip2(n11566), .s(n11472), .op(
        n6403) );
  mux2_1 U12638 ( .ip1(\cache_data[3][45] ), .ip2(n11567), .s(n11472), .op(
        n6402) );
  mux2_1 U12639 ( .ip1(\cache_data[3][46] ), .ip2(n11568), .s(n11472), .op(
        n6401) );
  mux2_1 U12640 ( .ip1(\cache_data[3][47] ), .ip2(n11569), .s(n11472), .op(
        n6400) );
  mux2_1 U12641 ( .ip1(\cache_data[3][48] ), .ip2(n11570), .s(n11472), .op(
        n6399) );
  mux2_1 U12642 ( .ip1(\cache_data[3][49] ), .ip2(n11571), .s(n11472), .op(
        n6398) );
  mux2_1 U12643 ( .ip1(\cache_data[3][50] ), .ip2(n11572), .s(n11472), .op(
        n6397) );
  buf_1 U12644 ( .ip(n11472), .op(n11473) );
  mux2_1 U12645 ( .ip1(\cache_data[3][51] ), .ip2(n11573), .s(n11473), .op(
        n6396) );
  mux2_1 U12646 ( .ip1(\cache_data[3][52] ), .ip2(n11574), .s(n11473), .op(
        n6395) );
  mux2_1 U12647 ( .ip1(\cache_data[3][53] ), .ip2(n11575), .s(n11473), .op(
        n6394) );
  mux2_1 U12648 ( .ip1(\cache_data[3][54] ), .ip2(n11576), .s(n11473), .op(
        n6393) );
  mux2_1 U12649 ( .ip1(\cache_data[3][55] ), .ip2(n11577), .s(n11473), .op(
        n6392) );
  mux2_1 U12650 ( .ip1(\cache_data[3][56] ), .ip2(n11578), .s(n11472), .op(
        n6391) );
  mux2_1 U12651 ( .ip1(\cache_data[3][57] ), .ip2(n11580), .s(n11472), .op(
        n6390) );
  mux2_1 U12652 ( .ip1(\cache_data[3][58] ), .ip2(n11581), .s(n11473), .op(
        n6389) );
  mux2_1 U12653 ( .ip1(\cache_data[3][59] ), .ip2(n11582), .s(n11473), .op(
        n6388) );
  mux2_1 U12654 ( .ip1(\cache_data[3][60] ), .ip2(n11583), .s(n11473), .op(
        n6387) );
  mux2_1 U12655 ( .ip1(\cache_data[3][61] ), .ip2(n11584), .s(n11473), .op(
        n6386) );
  mux2_1 U12656 ( .ip1(\cache_data[3][62] ), .ip2(n11585), .s(n11473), .op(
        n6385) );
  mux2_1 U12657 ( .ip1(\cache_data[3][63] ), .ip2(n11587), .s(n11473), .op(
        n6384) );
  nor2_1 U12658 ( .ip1(n11609), .ip2(n11476), .op(n11474) );
  mux2_1 U12659 ( .ip1(\cache_data[3][64] ), .ip2(n11554), .s(n11474), .op(
        n6383) );
  mux2_1 U12660 ( .ip1(\cache_data[3][65] ), .ip2(n11555), .s(n11474), .op(
        n6382) );
  mux2_1 U12661 ( .ip1(\cache_data[3][66] ), .ip2(n11556), .s(n11474), .op(
        n6381) );
  mux2_1 U12662 ( .ip1(\cache_data[3][67] ), .ip2(n11557), .s(n11474), .op(
        n6380) );
  mux2_1 U12663 ( .ip1(\cache_data[3][68] ), .ip2(n11558), .s(n11474), .op(
        n6379) );
  mux2_1 U12664 ( .ip1(\cache_data[3][69] ), .ip2(n11559), .s(n11474), .op(
        n6378) );
  mux2_1 U12665 ( .ip1(\cache_data[3][70] ), .ip2(n11560), .s(n11474), .op(
        n6377) );
  mux2_1 U12666 ( .ip1(\cache_data[3][71] ), .ip2(n11561), .s(n11474), .op(
        n6376) );
  mux2_1 U12667 ( .ip1(\cache_data[3][72] ), .ip2(n11562), .s(n11474), .op(
        n6375) );
  mux2_1 U12668 ( .ip1(\cache_data[3][73] ), .ip2(n11563), .s(n11474), .op(
        n6374) );
  mux2_1 U12669 ( .ip1(\cache_data[3][74] ), .ip2(n11564), .s(n11474), .op(
        n6373) );
  mux2_1 U12670 ( .ip1(\cache_data[3][75] ), .ip2(n11565), .s(n11474), .op(
        n6372) );
  mux2_1 U12671 ( .ip1(\cache_data[3][76] ), .ip2(n11566), .s(n11474), .op(
        n6371) );
  mux2_1 U12672 ( .ip1(\cache_data[3][77] ), .ip2(n11567), .s(n11474), .op(
        n6370) );
  mux2_1 U12673 ( .ip1(\cache_data[3][78] ), .ip2(n11568), .s(n11474), .op(
        n6369) );
  mux2_1 U12674 ( .ip1(\cache_data[3][79] ), .ip2(n11569), .s(n11474), .op(
        n6368) );
  mux2_1 U12675 ( .ip1(\cache_data[3][80] ), .ip2(n11570), .s(n11474), .op(
        n6367) );
  mux2_1 U12676 ( .ip1(\cache_data[3][81] ), .ip2(n11571), .s(n11474), .op(
        n6366) );
  mux2_1 U12677 ( .ip1(\cache_data[3][82] ), .ip2(n11572), .s(n11474), .op(
        n6365) );
  buf_1 U12678 ( .ip(n11474), .op(n11475) );
  mux2_1 U12679 ( .ip1(\cache_data[3][83] ), .ip2(n11573), .s(n11475), .op(
        n6364) );
  mux2_1 U12680 ( .ip1(\cache_data[3][84] ), .ip2(n11574), .s(n11475), .op(
        n6363) );
  mux2_1 U12681 ( .ip1(\cache_data[3][85] ), .ip2(n11575), .s(n11475), .op(
        n6362) );
  mux2_1 U12682 ( .ip1(\cache_data[3][86] ), .ip2(n11576), .s(n11475), .op(
        n6361) );
  mux2_1 U12683 ( .ip1(\cache_data[3][87] ), .ip2(n11577), .s(n11475), .op(
        n6360) );
  mux2_1 U12684 ( .ip1(\cache_data[3][88] ), .ip2(n11578), .s(n11474), .op(
        n6359) );
  mux2_1 U12685 ( .ip1(\cache_data[3][89] ), .ip2(n11580), .s(n11474), .op(
        n6358) );
  mux2_1 U12686 ( .ip1(\cache_data[3][90] ), .ip2(n11581), .s(n11475), .op(
        n6357) );
  mux2_1 U12687 ( .ip1(\cache_data[3][91] ), .ip2(n11582), .s(n11475), .op(
        n6356) );
  mux2_1 U12688 ( .ip1(\cache_data[3][92] ), .ip2(n11583), .s(n11475), .op(
        n6355) );
  mux2_1 U12689 ( .ip1(\cache_data[3][93] ), .ip2(n11584), .s(n11475), .op(
        n6354) );
  mux2_1 U12690 ( .ip1(\cache_data[3][94] ), .ip2(n11585), .s(n11475), .op(
        n6353) );
  mux2_1 U12691 ( .ip1(\cache_data[3][95] ), .ip2(n11587), .s(n11475), .op(
        n6352) );
  nor2_1 U12692 ( .ip1(n11613), .ip2(n11476), .op(n11477) );
  mux2_1 U12693 ( .ip1(\cache_data[3][96] ), .ip2(n11554), .s(n11477), .op(
        n6351) );
  mux2_1 U12694 ( .ip1(\cache_data[3][97] ), .ip2(n11555), .s(n11477), .op(
        n6350) );
  mux2_1 U12695 ( .ip1(\cache_data[3][98] ), .ip2(n11556), .s(n11477), .op(
        n6349) );
  mux2_1 U12696 ( .ip1(\cache_data[3][99] ), .ip2(n11557), .s(n11477), .op(
        n6348) );
  mux2_1 U12697 ( .ip1(\cache_data[3][100] ), .ip2(n11558), .s(n11477), .op(
        n6347) );
  mux2_1 U12698 ( .ip1(\cache_data[3][101] ), .ip2(n11559), .s(n11477), .op(
        n6346) );
  mux2_1 U12699 ( .ip1(\cache_data[3][102] ), .ip2(n11560), .s(n11477), .op(
        n6345) );
  mux2_1 U12700 ( .ip1(\cache_data[3][103] ), .ip2(n11561), .s(n11477), .op(
        n6344) );
  mux2_1 U12701 ( .ip1(\cache_data[3][104] ), .ip2(n11562), .s(n11477), .op(
        n6343) );
  mux2_1 U12702 ( .ip1(\cache_data[3][105] ), .ip2(n11563), .s(n11477), .op(
        n6342) );
  mux2_1 U12703 ( .ip1(\cache_data[3][106] ), .ip2(n11564), .s(n11477), .op(
        n6341) );
  mux2_1 U12704 ( .ip1(\cache_data[3][107] ), .ip2(n11565), .s(n11477), .op(
        n6340) );
  mux2_1 U12705 ( .ip1(\cache_data[3][108] ), .ip2(n11566), .s(n11477), .op(
        n6339) );
  mux2_1 U12706 ( .ip1(\cache_data[3][109] ), .ip2(n11567), .s(n11477), .op(
        n6338) );
  mux2_1 U12707 ( .ip1(\cache_data[3][110] ), .ip2(n11568), .s(n11477), .op(
        n6337) );
  mux2_1 U12708 ( .ip1(\cache_data[3][111] ), .ip2(n11569), .s(n11477), .op(
        n6336) );
  mux2_1 U12709 ( .ip1(\cache_data[3][112] ), .ip2(n11570), .s(n11477), .op(
        n6335) );
  mux2_1 U12710 ( .ip1(\cache_data[3][113] ), .ip2(n11571), .s(n11477), .op(
        n6334) );
  mux2_1 U12711 ( .ip1(\cache_data[3][114] ), .ip2(n11572), .s(n11477), .op(
        n6333) );
  buf_1 U12712 ( .ip(n11477), .op(n11478) );
  mux2_1 U12713 ( .ip1(\cache_data[3][115] ), .ip2(n11573), .s(n11478), .op(
        n6332) );
  mux2_1 U12714 ( .ip1(\cache_data[3][116] ), .ip2(n11574), .s(n11478), .op(
        n6331) );
  mux2_1 U12715 ( .ip1(\cache_data[3][117] ), .ip2(n11575), .s(n11478), .op(
        n6330) );
  mux2_1 U12716 ( .ip1(\cache_data[3][118] ), .ip2(n11576), .s(n11478), .op(
        n6329) );
  mux2_1 U12717 ( .ip1(\cache_data[3][119] ), .ip2(n11577), .s(n11478), .op(
        n6328) );
  mux2_1 U12718 ( .ip1(\cache_data[3][120] ), .ip2(n11578), .s(n11477), .op(
        n6327) );
  mux2_1 U12719 ( .ip1(\cache_data[3][121] ), .ip2(n11580), .s(n11477), .op(
        n6326) );
  mux2_1 U12720 ( .ip1(\cache_data[3][122] ), .ip2(n11581), .s(n11478), .op(
        n6325) );
  mux2_1 U12721 ( .ip1(\cache_data[3][123] ), .ip2(n11582), .s(n11478), .op(
        n6324) );
  mux2_1 U12722 ( .ip1(\cache_data[3][124] ), .ip2(n11583), .s(n11478), .op(
        n6323) );
  mux2_1 U12723 ( .ip1(\cache_data[3][125] ), .ip2(n11584), .s(n11478), .op(
        n6322) );
  mux2_1 U12724 ( .ip1(\cache_data[3][126] ), .ip2(n11585), .s(n11478), .op(
        n6321) );
  mux2_1 U12725 ( .ip1(\cache_data[3][127] ), .ip2(n11587), .s(n11478), .op(
        n6320) );
  nor2_1 U12726 ( .ip1(n11603), .ip2(n8136), .op(n11479) );
  mux2_1 U12727 ( .ip1(\cache_data[4][0] ), .ip2(n11554), .s(n11479), .op(
        n6319) );
  mux2_1 U12728 ( .ip1(\cache_data[4][1] ), .ip2(n11555), .s(n11479), .op(
        n6318) );
  mux2_1 U12729 ( .ip1(\cache_data[4][2] ), .ip2(n11556), .s(n11479), .op(
        n6317) );
  mux2_1 U12730 ( .ip1(\cache_data[4][3] ), .ip2(n11557), .s(n11479), .op(
        n6316) );
  mux2_1 U12731 ( .ip1(\cache_data[4][4] ), .ip2(n11558), .s(n11479), .op(
        n6315) );
  mux2_1 U12732 ( .ip1(\cache_data[4][5] ), .ip2(n11559), .s(n11479), .op(
        n6314) );
  mux2_1 U12733 ( .ip1(\cache_data[4][6] ), .ip2(n11560), .s(n11479), .op(
        n6313) );
  mux2_1 U12734 ( .ip1(\cache_data[4][7] ), .ip2(n11561), .s(n11479), .op(
        n6312) );
  mux2_1 U12735 ( .ip1(\cache_data[4][8] ), .ip2(n11562), .s(n11479), .op(
        n6311) );
  mux2_1 U12736 ( .ip1(\cache_data[4][9] ), .ip2(n11563), .s(n11479), .op(
        n6310) );
  mux2_1 U12737 ( .ip1(\cache_data[4][10] ), .ip2(n11564), .s(n11479), .op(
        n6309) );
  mux2_1 U12738 ( .ip1(\cache_data[4][11] ), .ip2(n11565), .s(n11479), .op(
        n6308) );
  mux2_1 U12739 ( .ip1(\cache_data[4][12] ), .ip2(n11566), .s(n11479), .op(
        n6307) );
  mux2_1 U12740 ( .ip1(\cache_data[4][13] ), .ip2(n11567), .s(n11479), .op(
        n6306) );
  mux2_1 U12741 ( .ip1(\cache_data[4][14] ), .ip2(n11568), .s(n11479), .op(
        n6305) );
  mux2_1 U12742 ( .ip1(\cache_data[4][15] ), .ip2(n11569), .s(n11479), .op(
        n6304) );
  mux2_1 U12743 ( .ip1(\cache_data[4][16] ), .ip2(n11570), .s(n11479), .op(
        n6303) );
  mux2_1 U12744 ( .ip1(\cache_data[4][17] ), .ip2(n11571), .s(n11479), .op(
        n6302) );
  mux2_1 U12745 ( .ip1(\cache_data[4][18] ), .ip2(n11572), .s(n11479), .op(
        n6301) );
  buf_1 U12746 ( .ip(n11479), .op(n11480) );
  mux2_1 U12747 ( .ip1(\cache_data[4][19] ), .ip2(n11573), .s(n11480), .op(
        n6300) );
  mux2_1 U12748 ( .ip1(\cache_data[4][20] ), .ip2(n11574), .s(n11480), .op(
        n6299) );
  mux2_1 U12749 ( .ip1(\cache_data[4][21] ), .ip2(n11575), .s(n11480), .op(
        n6298) );
  mux2_1 U12750 ( .ip1(\cache_data[4][22] ), .ip2(n11576), .s(n11480), .op(
        n6297) );
  mux2_1 U12751 ( .ip1(\cache_data[4][23] ), .ip2(n11577), .s(n11480), .op(
        n6296) );
  mux2_1 U12752 ( .ip1(\cache_data[4][24] ), .ip2(n11578), .s(n11479), .op(
        n6295) );
  mux2_1 U12753 ( .ip1(\cache_data[4][25] ), .ip2(n11580), .s(n11479), .op(
        n6294) );
  mux2_1 U12754 ( .ip1(\cache_data[4][26] ), .ip2(n11581), .s(n11480), .op(
        n6293) );
  mux2_1 U12755 ( .ip1(\cache_data[4][27] ), .ip2(n11582), .s(n11480), .op(
        n6292) );
  mux2_1 U12756 ( .ip1(\cache_data[4][28] ), .ip2(n11583), .s(n11480), .op(
        n6291) );
  mux2_1 U12757 ( .ip1(\cache_data[4][29] ), .ip2(n11584), .s(n11480), .op(
        n6290) );
  mux2_1 U12758 ( .ip1(\cache_data[4][30] ), .ip2(n11585), .s(n11480), .op(
        n6289) );
  mux2_1 U12759 ( .ip1(\cache_data[4][31] ), .ip2(n11587), .s(n11480), .op(
        n6288) );
  nor2_1 U12760 ( .ip1(n11606), .ip2(n8136), .op(n11481) );
  mux2_1 U12761 ( .ip1(\cache_data[4][32] ), .ip2(n11554), .s(n11481), .op(
        n6287) );
  mux2_1 U12762 ( .ip1(\cache_data[4][33] ), .ip2(n11555), .s(n11481), .op(
        n6286) );
  mux2_1 U12763 ( .ip1(\cache_data[4][34] ), .ip2(n11556), .s(n11481), .op(
        n6285) );
  mux2_1 U12764 ( .ip1(\cache_data[4][35] ), .ip2(n11557), .s(n11481), .op(
        n6284) );
  mux2_1 U12765 ( .ip1(\cache_data[4][36] ), .ip2(n11558), .s(n11481), .op(
        n6283) );
  mux2_1 U12766 ( .ip1(\cache_data[4][37] ), .ip2(n11559), .s(n11481), .op(
        n6282) );
  mux2_1 U12767 ( .ip1(\cache_data[4][38] ), .ip2(n11560), .s(n11481), .op(
        n6281) );
  mux2_1 U12768 ( .ip1(\cache_data[4][39] ), .ip2(n11561), .s(n11481), .op(
        n6280) );
  mux2_1 U12769 ( .ip1(\cache_data[4][40] ), .ip2(n11562), .s(n11481), .op(
        n6279) );
  mux2_1 U12770 ( .ip1(\cache_data[4][41] ), .ip2(n11563), .s(n11481), .op(
        n6278) );
  mux2_1 U12771 ( .ip1(\cache_data[4][42] ), .ip2(n11564), .s(n11481), .op(
        n6277) );
  mux2_1 U12772 ( .ip1(\cache_data[4][43] ), .ip2(n11565), .s(n11481), .op(
        n6276) );
  mux2_1 U12773 ( .ip1(\cache_data[4][44] ), .ip2(n11566), .s(n11481), .op(
        n6275) );
  mux2_1 U12774 ( .ip1(\cache_data[4][45] ), .ip2(n11567), .s(n11481), .op(
        n6274) );
  mux2_1 U12775 ( .ip1(\cache_data[4][46] ), .ip2(n11568), .s(n11481), .op(
        n6273) );
  mux2_1 U12776 ( .ip1(\cache_data[4][47] ), .ip2(n11569), .s(n11481), .op(
        n6272) );
  mux2_1 U12777 ( .ip1(\cache_data[4][48] ), .ip2(n11570), .s(n11481), .op(
        n6271) );
  mux2_1 U12778 ( .ip1(\cache_data[4][49] ), .ip2(n11571), .s(n11481), .op(
        n6270) );
  mux2_1 U12779 ( .ip1(\cache_data[4][50] ), .ip2(n11572), .s(n11481), .op(
        n6269) );
  buf_1 U12780 ( .ip(n11481), .op(n11482) );
  mux2_1 U12781 ( .ip1(\cache_data[4][51] ), .ip2(n11573), .s(n11482), .op(
        n6268) );
  mux2_1 U12782 ( .ip1(\cache_data[4][52] ), .ip2(n11574), .s(n11482), .op(
        n6267) );
  mux2_1 U12783 ( .ip1(\cache_data[4][53] ), .ip2(n11575), .s(n11482), .op(
        n6266) );
  mux2_1 U12784 ( .ip1(\cache_data[4][54] ), .ip2(n11576), .s(n11482), .op(
        n6265) );
  mux2_1 U12785 ( .ip1(\cache_data[4][55] ), .ip2(n11577), .s(n11482), .op(
        n6264) );
  mux2_1 U12786 ( .ip1(\cache_data[4][56] ), .ip2(n11578), .s(n11481), .op(
        n6263) );
  mux2_1 U12787 ( .ip1(\cache_data[4][57] ), .ip2(n11580), .s(n11481), .op(
        n6262) );
  mux2_1 U12788 ( .ip1(\cache_data[4][58] ), .ip2(n11581), .s(n11482), .op(
        n6261) );
  mux2_1 U12789 ( .ip1(\cache_data[4][59] ), .ip2(n11582), .s(n11482), .op(
        n6260) );
  mux2_1 U12790 ( .ip1(\cache_data[4][60] ), .ip2(n11583), .s(n11482), .op(
        n6259) );
  mux2_1 U12791 ( .ip1(\cache_data[4][61] ), .ip2(n11584), .s(n11482), .op(
        n6258) );
  mux2_1 U12792 ( .ip1(\cache_data[4][62] ), .ip2(n11585), .s(n11482), .op(
        n6257) );
  mux2_1 U12793 ( .ip1(\cache_data[4][63] ), .ip2(n11587), .s(n11482), .op(
        n6256) );
  nor2_1 U12794 ( .ip1(n11609), .ip2(n8136), .op(n11483) );
  mux2_1 U12795 ( .ip1(\cache_data[4][64] ), .ip2(n11554), .s(n11483), .op(
        n6255) );
  mux2_1 U12796 ( .ip1(\cache_data[4][65] ), .ip2(n11555), .s(n11483), .op(
        n6254) );
  mux2_1 U12797 ( .ip1(\cache_data[4][66] ), .ip2(n11556), .s(n11483), .op(
        n6253) );
  mux2_1 U12798 ( .ip1(\cache_data[4][67] ), .ip2(n11557), .s(n11483), .op(
        n6252) );
  mux2_1 U12799 ( .ip1(\cache_data[4][68] ), .ip2(n11558), .s(n11483), .op(
        n6251) );
  mux2_1 U12800 ( .ip1(\cache_data[4][69] ), .ip2(n11559), .s(n11483), .op(
        n6250) );
  mux2_1 U12801 ( .ip1(\cache_data[4][70] ), .ip2(n11560), .s(n11483), .op(
        n6249) );
  mux2_1 U12802 ( .ip1(\cache_data[4][71] ), .ip2(n11561), .s(n11483), .op(
        n6248) );
  mux2_1 U12803 ( .ip1(\cache_data[4][72] ), .ip2(n11562), .s(n11483), .op(
        n6247) );
  mux2_1 U12804 ( .ip1(\cache_data[4][73] ), .ip2(n11563), .s(n11483), .op(
        n6246) );
  mux2_1 U12805 ( .ip1(\cache_data[4][74] ), .ip2(n11564), .s(n11483), .op(
        n6245) );
  mux2_1 U12806 ( .ip1(\cache_data[4][75] ), .ip2(n11565), .s(n11483), .op(
        n6244) );
  mux2_1 U12807 ( .ip1(\cache_data[4][76] ), .ip2(n11566), .s(n11483), .op(
        n6243) );
  mux2_1 U12808 ( .ip1(\cache_data[4][77] ), .ip2(n11567), .s(n11483), .op(
        n6242) );
  mux2_1 U12809 ( .ip1(\cache_data[4][78] ), .ip2(n11568), .s(n11483), .op(
        n6241) );
  mux2_1 U12810 ( .ip1(\cache_data[4][79] ), .ip2(n11569), .s(n11483), .op(
        n6240) );
  mux2_1 U12811 ( .ip1(\cache_data[4][80] ), .ip2(n11570), .s(n11483), .op(
        n6239) );
  mux2_1 U12812 ( .ip1(\cache_data[4][81] ), .ip2(n11571), .s(n11483), .op(
        n6238) );
  mux2_1 U12813 ( .ip1(\cache_data[4][82] ), .ip2(n11572), .s(n11483), .op(
        n6237) );
  buf_1 U12814 ( .ip(n11483), .op(n11484) );
  mux2_1 U12815 ( .ip1(\cache_data[4][83] ), .ip2(n11573), .s(n11484), .op(
        n6236) );
  mux2_1 U12816 ( .ip1(\cache_data[4][84] ), .ip2(n11574), .s(n11484), .op(
        n6235) );
  mux2_1 U12817 ( .ip1(\cache_data[4][85] ), .ip2(n11575), .s(n11484), .op(
        n6234) );
  mux2_1 U12818 ( .ip1(\cache_data[4][86] ), .ip2(n11576), .s(n11484), .op(
        n6233) );
  mux2_1 U12819 ( .ip1(\cache_data[4][87] ), .ip2(n11577), .s(n11484), .op(
        n6232) );
  mux2_1 U12820 ( .ip1(\cache_data[4][88] ), .ip2(n11578), .s(n11483), .op(
        n6231) );
  mux2_1 U12821 ( .ip1(\cache_data[4][89] ), .ip2(n11580), .s(n11483), .op(
        n6230) );
  mux2_1 U12822 ( .ip1(\cache_data[4][90] ), .ip2(n11581), .s(n11484), .op(
        n6229) );
  mux2_1 U12823 ( .ip1(\cache_data[4][91] ), .ip2(n11582), .s(n11484), .op(
        n6228) );
  mux2_1 U12824 ( .ip1(\cache_data[4][92] ), .ip2(n11583), .s(n11484), .op(
        n6227) );
  mux2_1 U12825 ( .ip1(\cache_data[4][93] ), .ip2(n11584), .s(n11484), .op(
        n6226) );
  mux2_1 U12826 ( .ip1(\cache_data[4][94] ), .ip2(n11585), .s(n11484), .op(
        n6225) );
  mux2_1 U12827 ( .ip1(\cache_data[4][95] ), .ip2(n11587), .s(n11484), .op(
        n6224) );
  nor2_1 U12828 ( .ip1(n11613), .ip2(n8136), .op(n11485) );
  mux2_1 U12829 ( .ip1(\cache_data[4][96] ), .ip2(n11554), .s(n11485), .op(
        n6223) );
  mux2_1 U12830 ( .ip1(\cache_data[4][97] ), .ip2(n11555), .s(n11485), .op(
        n6222) );
  mux2_1 U12831 ( .ip1(\cache_data[4][98] ), .ip2(n11556), .s(n11485), .op(
        n6221) );
  mux2_1 U12832 ( .ip1(\cache_data[4][99] ), .ip2(n11557), .s(n11485), .op(
        n6220) );
  mux2_1 U12833 ( .ip1(\cache_data[4][100] ), .ip2(n11558), .s(n11485), .op(
        n6219) );
  mux2_1 U12834 ( .ip1(\cache_data[4][101] ), .ip2(n11559), .s(n11485), .op(
        n6218) );
  mux2_1 U12835 ( .ip1(\cache_data[4][102] ), .ip2(n11560), .s(n11485), .op(
        n6217) );
  mux2_1 U12836 ( .ip1(\cache_data[4][103] ), .ip2(n11561), .s(n11485), .op(
        n6216) );
  mux2_1 U12837 ( .ip1(\cache_data[4][104] ), .ip2(n11562), .s(n11485), .op(
        n6215) );
  mux2_1 U12838 ( .ip1(\cache_data[4][105] ), .ip2(n11563), .s(n11485), .op(
        n6214) );
  mux2_1 U12839 ( .ip1(\cache_data[4][106] ), .ip2(n11564), .s(n11485), .op(
        n6213) );
  mux2_1 U12840 ( .ip1(\cache_data[4][107] ), .ip2(n11565), .s(n11485), .op(
        n6212) );
  mux2_1 U12841 ( .ip1(\cache_data[4][108] ), .ip2(n11566), .s(n11485), .op(
        n6211) );
  mux2_1 U12842 ( .ip1(\cache_data[4][109] ), .ip2(n11567), .s(n11485), .op(
        n6210) );
  mux2_1 U12843 ( .ip1(\cache_data[4][110] ), .ip2(n11568), .s(n11485), .op(
        n6209) );
  mux2_1 U12844 ( .ip1(\cache_data[4][111] ), .ip2(n11569), .s(n11485), .op(
        n6208) );
  mux2_1 U12845 ( .ip1(\cache_data[4][112] ), .ip2(n11570), .s(n11485), .op(
        n6207) );
  mux2_1 U12846 ( .ip1(\cache_data[4][113] ), .ip2(n11571), .s(n11485), .op(
        n6206) );
  mux2_1 U12847 ( .ip1(\cache_data[4][114] ), .ip2(n11572), .s(n11485), .op(
        n6205) );
  buf_1 U12848 ( .ip(n11485), .op(n11486) );
  mux2_1 U12849 ( .ip1(\cache_data[4][115] ), .ip2(n11573), .s(n11486), .op(
        n6204) );
  mux2_1 U12850 ( .ip1(\cache_data[4][116] ), .ip2(n11574), .s(n11486), .op(
        n6203) );
  mux2_1 U12851 ( .ip1(\cache_data[4][117] ), .ip2(n11575), .s(n11486), .op(
        n6202) );
  mux2_1 U12852 ( .ip1(\cache_data[4][118] ), .ip2(n11576), .s(n11486), .op(
        n6201) );
  mux2_1 U12853 ( .ip1(\cache_data[4][119] ), .ip2(n11577), .s(n11486), .op(
        n6200) );
  mux2_1 U12854 ( .ip1(\cache_data[4][120] ), .ip2(n11578), .s(n11485), .op(
        n6199) );
  mux2_1 U12855 ( .ip1(\cache_data[4][121] ), .ip2(n11580), .s(n11485), .op(
        n6198) );
  mux2_1 U12856 ( .ip1(\cache_data[4][122] ), .ip2(n11581), .s(n11486), .op(
        n6197) );
  mux2_1 U12857 ( .ip1(\cache_data[4][123] ), .ip2(n11582), .s(n11486), .op(
        n6196) );
  mux2_1 U12858 ( .ip1(\cache_data[4][124] ), .ip2(n11583), .s(n11486), .op(
        n6195) );
  mux2_1 U12859 ( .ip1(\cache_data[4][125] ), .ip2(n11584), .s(n11486), .op(
        n6194) );
  mux2_1 U12860 ( .ip1(\cache_data[4][126] ), .ip2(n11585), .s(n11486), .op(
        n6193) );
  mux2_1 U12861 ( .ip1(\cache_data[4][127] ), .ip2(n11587), .s(n11486), .op(
        n6192) );
  nor2_1 U12862 ( .ip1(n11603), .ip2(n11493), .op(n11487) );
  mux2_1 U12863 ( .ip1(\cache_data[5][0] ), .ip2(n11554), .s(n11487), .op(
        n6191) );
  mux2_1 U12864 ( .ip1(\cache_data[5][1] ), .ip2(n11555), .s(n11487), .op(
        n6190) );
  mux2_1 U12865 ( .ip1(\cache_data[5][2] ), .ip2(n11556), .s(n11487), .op(
        n6189) );
  mux2_1 U12866 ( .ip1(\cache_data[5][3] ), .ip2(n11557), .s(n11487), .op(
        n6188) );
  mux2_1 U12867 ( .ip1(\cache_data[5][4] ), .ip2(n11558), .s(n11487), .op(
        n6187) );
  mux2_1 U12868 ( .ip1(\cache_data[5][5] ), .ip2(n11559), .s(n11487), .op(
        n6186) );
  mux2_1 U12869 ( .ip1(\cache_data[5][6] ), .ip2(n11560), .s(n11487), .op(
        n6185) );
  mux2_1 U12870 ( .ip1(\cache_data[5][7] ), .ip2(n11561), .s(n11487), .op(
        n6184) );
  mux2_1 U12871 ( .ip1(\cache_data[5][8] ), .ip2(n11562), .s(n11487), .op(
        n6183) );
  mux2_1 U12872 ( .ip1(\cache_data[5][9] ), .ip2(n11563), .s(n11487), .op(
        n6182) );
  mux2_1 U12873 ( .ip1(\cache_data[5][10] ), .ip2(n11564), .s(n11487), .op(
        n6181) );
  mux2_1 U12874 ( .ip1(\cache_data[5][11] ), .ip2(n11565), .s(n11487), .op(
        n6180) );
  mux2_1 U12875 ( .ip1(\cache_data[5][12] ), .ip2(n11566), .s(n11487), .op(
        n6179) );
  mux2_1 U12876 ( .ip1(\cache_data[5][13] ), .ip2(n11567), .s(n11487), .op(
        n6178) );
  mux2_1 U12877 ( .ip1(\cache_data[5][14] ), .ip2(n11568), .s(n11487), .op(
        n6177) );
  mux2_1 U12878 ( .ip1(\cache_data[5][15] ), .ip2(n11569), .s(n11487), .op(
        n6176) );
  mux2_1 U12879 ( .ip1(\cache_data[5][16] ), .ip2(n11570), .s(n11487), .op(
        n6175) );
  mux2_1 U12880 ( .ip1(\cache_data[5][17] ), .ip2(n11571), .s(n11487), .op(
        n6174) );
  mux2_1 U12881 ( .ip1(\cache_data[5][18] ), .ip2(n11572), .s(n11487), .op(
        n6173) );
  buf_1 U12882 ( .ip(n11487), .op(n11488) );
  mux2_1 U12883 ( .ip1(\cache_data[5][19] ), .ip2(n11573), .s(n11488), .op(
        n6172) );
  mux2_1 U12884 ( .ip1(\cache_data[5][20] ), .ip2(n11574), .s(n11488), .op(
        n6171) );
  mux2_1 U12885 ( .ip1(\cache_data[5][21] ), .ip2(n11575), .s(n11488), .op(
        n6170) );
  mux2_1 U12886 ( .ip1(\cache_data[5][22] ), .ip2(n11576), .s(n11488), .op(
        n6169) );
  mux2_1 U12887 ( .ip1(\cache_data[5][23] ), .ip2(n11577), .s(n11488), .op(
        n6168) );
  mux2_1 U12888 ( .ip1(\cache_data[5][24] ), .ip2(n11578), .s(n11487), .op(
        n6167) );
  mux2_1 U12889 ( .ip1(\cache_data[5][25] ), .ip2(n11580), .s(n11487), .op(
        n6166) );
  mux2_1 U12890 ( .ip1(\cache_data[5][26] ), .ip2(n11581), .s(n11488), .op(
        n6165) );
  mux2_1 U12891 ( .ip1(\cache_data[5][27] ), .ip2(n11582), .s(n11488), .op(
        n6164) );
  mux2_1 U12892 ( .ip1(\cache_data[5][28] ), .ip2(n11583), .s(n11488), .op(
        n6163) );
  mux2_1 U12893 ( .ip1(\cache_data[5][29] ), .ip2(n11584), .s(n11488), .op(
        n6162) );
  mux2_1 U12894 ( .ip1(\cache_data[5][30] ), .ip2(n11585), .s(n11488), .op(
        n6161) );
  mux2_1 U12895 ( .ip1(\cache_data[5][31] ), .ip2(n11587), .s(n11488), .op(
        n6160) );
  nor2_1 U12896 ( .ip1(n11606), .ip2(n11493), .op(n11489) );
  mux2_1 U12897 ( .ip1(\cache_data[5][32] ), .ip2(n11554), .s(n11489), .op(
        n6159) );
  mux2_1 U12898 ( .ip1(\cache_data[5][33] ), .ip2(n11555), .s(n11489), .op(
        n6158) );
  mux2_1 U12899 ( .ip1(\cache_data[5][34] ), .ip2(n11556), .s(n11489), .op(
        n6157) );
  mux2_1 U12900 ( .ip1(\cache_data[5][35] ), .ip2(n11557), .s(n11489), .op(
        n6156) );
  mux2_1 U12901 ( .ip1(\cache_data[5][36] ), .ip2(n11558), .s(n11489), .op(
        n6155) );
  mux2_1 U12902 ( .ip1(\cache_data[5][37] ), .ip2(n11559), .s(n11489), .op(
        n6154) );
  mux2_1 U12903 ( .ip1(\cache_data[5][38] ), .ip2(n11560), .s(n11489), .op(
        n6153) );
  mux2_1 U12904 ( .ip1(\cache_data[5][39] ), .ip2(n11561), .s(n11489), .op(
        n6152) );
  mux2_1 U12905 ( .ip1(\cache_data[5][40] ), .ip2(n11562), .s(n11489), .op(
        n6151) );
  mux2_1 U12906 ( .ip1(\cache_data[5][41] ), .ip2(n11563), .s(n11489), .op(
        n6150) );
  mux2_1 U12907 ( .ip1(\cache_data[5][42] ), .ip2(n11564), .s(n11489), .op(
        n6149) );
  mux2_1 U12908 ( .ip1(\cache_data[5][43] ), .ip2(n11565), .s(n11489), .op(
        n6148) );
  mux2_1 U12909 ( .ip1(\cache_data[5][44] ), .ip2(n11566), .s(n11489), .op(
        n6147) );
  mux2_1 U12910 ( .ip1(\cache_data[5][45] ), .ip2(n11567), .s(n11489), .op(
        n6146) );
  mux2_1 U12911 ( .ip1(\cache_data[5][46] ), .ip2(n11568), .s(n11489), .op(
        n6145) );
  mux2_1 U12912 ( .ip1(\cache_data[5][47] ), .ip2(n11569), .s(n11489), .op(
        n6144) );
  mux2_1 U12913 ( .ip1(\cache_data[5][48] ), .ip2(n11570), .s(n11489), .op(
        n6143) );
  mux2_1 U12914 ( .ip1(\cache_data[5][49] ), .ip2(n11571), .s(n11489), .op(
        n6142) );
  mux2_1 U12915 ( .ip1(\cache_data[5][50] ), .ip2(n11572), .s(n11489), .op(
        n6141) );
  buf_1 U12916 ( .ip(n11489), .op(n11490) );
  mux2_1 U12917 ( .ip1(\cache_data[5][51] ), .ip2(n11573), .s(n11490), .op(
        n6140) );
  mux2_1 U12918 ( .ip1(\cache_data[5][52] ), .ip2(n11574), .s(n11490), .op(
        n6139) );
  mux2_1 U12919 ( .ip1(\cache_data[5][53] ), .ip2(n11575), .s(n11490), .op(
        n6138) );
  mux2_1 U12920 ( .ip1(\cache_data[5][54] ), .ip2(n11576), .s(n11490), .op(
        n6137) );
  mux2_1 U12921 ( .ip1(\cache_data[5][55] ), .ip2(n11577), .s(n11490), .op(
        n6136) );
  mux2_1 U12922 ( .ip1(\cache_data[5][56] ), .ip2(n11578), .s(n11489), .op(
        n6135) );
  mux2_1 U12923 ( .ip1(\cache_data[5][57] ), .ip2(n11580), .s(n11489), .op(
        n6134) );
  mux2_1 U12924 ( .ip1(\cache_data[5][58] ), .ip2(n11581), .s(n11490), .op(
        n6133) );
  mux2_1 U12925 ( .ip1(\cache_data[5][59] ), .ip2(n11582), .s(n11490), .op(
        n6132) );
  mux2_1 U12926 ( .ip1(\cache_data[5][60] ), .ip2(n11583), .s(n11490), .op(
        n6131) );
  mux2_1 U12927 ( .ip1(\cache_data[5][61] ), .ip2(n11584), .s(n11490), .op(
        n6130) );
  mux2_1 U12928 ( .ip1(\cache_data[5][62] ), .ip2(n11585), .s(n11490), .op(
        n6129) );
  mux2_1 U12929 ( .ip1(\cache_data[5][63] ), .ip2(n11587), .s(n11490), .op(
        n6128) );
  nor2_1 U12930 ( .ip1(n11609), .ip2(n11493), .op(n11491) );
  mux2_1 U12931 ( .ip1(\cache_data[5][64] ), .ip2(n11554), .s(n11491), .op(
        n6127) );
  mux2_1 U12932 ( .ip1(\cache_data[5][65] ), .ip2(n11555), .s(n11491), .op(
        n6126) );
  mux2_1 U12933 ( .ip1(\cache_data[5][66] ), .ip2(n11556), .s(n11491), .op(
        n6125) );
  mux2_1 U12934 ( .ip1(\cache_data[5][67] ), .ip2(n11557), .s(n11491), .op(
        n6124) );
  mux2_1 U12935 ( .ip1(\cache_data[5][68] ), .ip2(n11558), .s(n11491), .op(
        n6123) );
  mux2_1 U12936 ( .ip1(\cache_data[5][69] ), .ip2(n11559), .s(n11491), .op(
        n6122) );
  mux2_1 U12937 ( .ip1(\cache_data[5][70] ), .ip2(n11560), .s(n11491), .op(
        n6121) );
  mux2_1 U12938 ( .ip1(\cache_data[5][71] ), .ip2(n11561), .s(n11491), .op(
        n6120) );
  mux2_1 U12939 ( .ip1(\cache_data[5][72] ), .ip2(n11562), .s(n11491), .op(
        n6119) );
  mux2_1 U12940 ( .ip1(\cache_data[5][73] ), .ip2(n11563), .s(n11491), .op(
        n6118) );
  mux2_1 U12941 ( .ip1(\cache_data[5][74] ), .ip2(n11564), .s(n11491), .op(
        n6117) );
  mux2_1 U12942 ( .ip1(\cache_data[5][75] ), .ip2(n11565), .s(n11491), .op(
        n6116) );
  mux2_1 U12943 ( .ip1(\cache_data[5][76] ), .ip2(n11566), .s(n11491), .op(
        n6115) );
  mux2_1 U12944 ( .ip1(\cache_data[5][77] ), .ip2(n11567), .s(n11491), .op(
        n6114) );
  mux2_1 U12945 ( .ip1(\cache_data[5][78] ), .ip2(n11568), .s(n11491), .op(
        n6113) );
  mux2_1 U12946 ( .ip1(\cache_data[5][79] ), .ip2(n11569), .s(n11491), .op(
        n6112) );
  mux2_1 U12947 ( .ip1(\cache_data[5][80] ), .ip2(n11570), .s(n11491), .op(
        n6111) );
  mux2_1 U12948 ( .ip1(\cache_data[5][81] ), .ip2(n11571), .s(n11491), .op(
        n6110) );
  mux2_1 U12949 ( .ip1(\cache_data[5][82] ), .ip2(n11572), .s(n11491), .op(
        n6109) );
  buf_1 U12950 ( .ip(n11491), .op(n11492) );
  mux2_1 U12951 ( .ip1(\cache_data[5][83] ), .ip2(n11573), .s(n11492), .op(
        n6108) );
  mux2_1 U12952 ( .ip1(\cache_data[5][84] ), .ip2(n11574), .s(n11492), .op(
        n6107) );
  mux2_1 U12953 ( .ip1(\cache_data[5][85] ), .ip2(n11575), .s(n11492), .op(
        n6106) );
  mux2_1 U12954 ( .ip1(\cache_data[5][86] ), .ip2(n11576), .s(n11492), .op(
        n6105) );
  mux2_1 U12955 ( .ip1(\cache_data[5][87] ), .ip2(n11577), .s(n11492), .op(
        n6104) );
  mux2_1 U12956 ( .ip1(\cache_data[5][88] ), .ip2(n11578), .s(n11491), .op(
        n6103) );
  mux2_1 U12957 ( .ip1(\cache_data[5][89] ), .ip2(n11580), .s(n11491), .op(
        n6102) );
  mux2_1 U12958 ( .ip1(\cache_data[5][90] ), .ip2(n11581), .s(n11492), .op(
        n6101) );
  mux2_1 U12959 ( .ip1(\cache_data[5][91] ), .ip2(n11582), .s(n11492), .op(
        n6100) );
  mux2_1 U12960 ( .ip1(\cache_data[5][92] ), .ip2(n11583), .s(n11492), .op(
        n6099) );
  mux2_1 U12961 ( .ip1(\cache_data[5][93] ), .ip2(n11584), .s(n11492), .op(
        n6098) );
  mux2_1 U12962 ( .ip1(\cache_data[5][94] ), .ip2(n11585), .s(n11492), .op(
        n6097) );
  mux2_1 U12963 ( .ip1(\cache_data[5][95] ), .ip2(n11587), .s(n11492), .op(
        n6096) );
  nor2_1 U12964 ( .ip1(n11613), .ip2(n11493), .op(n11494) );
  mux2_1 U12965 ( .ip1(\cache_data[5][96] ), .ip2(n11554), .s(n11494), .op(
        n6095) );
  mux2_1 U12966 ( .ip1(\cache_data[5][97] ), .ip2(n11555), .s(n11494), .op(
        n6094) );
  mux2_1 U12967 ( .ip1(\cache_data[5][98] ), .ip2(n11556), .s(n11494), .op(
        n6093) );
  mux2_1 U12968 ( .ip1(\cache_data[5][99] ), .ip2(n11557), .s(n11494), .op(
        n6092) );
  mux2_1 U12969 ( .ip1(\cache_data[5][100] ), .ip2(n11558), .s(n11494), .op(
        n6091) );
  mux2_1 U12970 ( .ip1(\cache_data[5][101] ), .ip2(n11559), .s(n11494), .op(
        n6090) );
  mux2_1 U12971 ( .ip1(\cache_data[5][102] ), .ip2(n11560), .s(n11494), .op(
        n6089) );
  mux2_1 U12972 ( .ip1(\cache_data[5][103] ), .ip2(n11561), .s(n11494), .op(
        n6088) );
  mux2_1 U12973 ( .ip1(\cache_data[5][104] ), .ip2(n11562), .s(n11494), .op(
        n6087) );
  mux2_1 U12974 ( .ip1(\cache_data[5][105] ), .ip2(n11563), .s(n11494), .op(
        n6086) );
  mux2_1 U12975 ( .ip1(\cache_data[5][106] ), .ip2(n11564), .s(n11494), .op(
        n6085) );
  mux2_1 U12976 ( .ip1(\cache_data[5][107] ), .ip2(n11565), .s(n11494), .op(
        n6084) );
  mux2_1 U12977 ( .ip1(\cache_data[5][108] ), .ip2(n11566), .s(n11494), .op(
        n6083) );
  mux2_1 U12978 ( .ip1(\cache_data[5][109] ), .ip2(n11567), .s(n11494), .op(
        n6082) );
  mux2_1 U12979 ( .ip1(\cache_data[5][110] ), .ip2(n11568), .s(n11494), .op(
        n6081) );
  mux2_1 U12980 ( .ip1(\cache_data[5][111] ), .ip2(n11569), .s(n11494), .op(
        n6080) );
  mux2_1 U12981 ( .ip1(\cache_data[5][112] ), .ip2(n11570), .s(n11494), .op(
        n6079) );
  mux2_1 U12982 ( .ip1(\cache_data[5][113] ), .ip2(n11571), .s(n11494), .op(
        n6078) );
  mux2_1 U12983 ( .ip1(\cache_data[5][114] ), .ip2(n11572), .s(n11494), .op(
        n6077) );
  buf_1 U12984 ( .ip(n11494), .op(n11495) );
  mux2_1 U12985 ( .ip1(\cache_data[5][115] ), .ip2(n11573), .s(n11495), .op(
        n6076) );
  mux2_1 U12986 ( .ip1(\cache_data[5][116] ), .ip2(n11574), .s(n11495), .op(
        n6075) );
  mux2_1 U12987 ( .ip1(\cache_data[5][117] ), .ip2(n11575), .s(n11495), .op(
        n6074) );
  mux2_1 U12988 ( .ip1(\cache_data[5][118] ), .ip2(n11576), .s(n11495), .op(
        n6073) );
  mux2_1 U12989 ( .ip1(\cache_data[5][119] ), .ip2(n11577), .s(n11495), .op(
        n6072) );
  mux2_1 U12990 ( .ip1(\cache_data[5][120] ), .ip2(n11578), .s(n11494), .op(
        n6071) );
  mux2_1 U12991 ( .ip1(\cache_data[5][121] ), .ip2(n11580), .s(n11494), .op(
        n6070) );
  mux2_1 U12992 ( .ip1(\cache_data[5][122] ), .ip2(n11581), .s(n11495), .op(
        n6069) );
  mux2_1 U12993 ( .ip1(\cache_data[5][123] ), .ip2(n11582), .s(n11495), .op(
        n6068) );
  mux2_1 U12994 ( .ip1(\cache_data[5][124] ), .ip2(n11583), .s(n11495), .op(
        n6067) );
  mux2_1 U12995 ( .ip1(\cache_data[5][125] ), .ip2(n11584), .s(n11495), .op(
        n6066) );
  mux2_1 U12996 ( .ip1(\cache_data[5][126] ), .ip2(n11585), .s(n11495), .op(
        n6065) );
  mux2_1 U12997 ( .ip1(\cache_data[5][127] ), .ip2(n11587), .s(n11495), .op(
        n6064) );
  buf_1 U12998 ( .ip(n11554), .op(n11614) );
  nor2_1 U12999 ( .ip1(n11603), .ip2(n11502), .op(n11496) );
  mux2_1 U13000 ( .ip1(\cache_data[6][0] ), .ip2(n11614), .s(n11496), .op(
        n6063) );
  buf_1 U13001 ( .ip(n11555), .op(n11615) );
  mux2_1 U13002 ( .ip1(\cache_data[6][1] ), .ip2(n11615), .s(n11496), .op(
        n6062) );
  buf_1 U13003 ( .ip(n11556), .op(n11616) );
  mux2_1 U13004 ( .ip1(\cache_data[6][2] ), .ip2(n11616), .s(n11496), .op(
        n6061) );
  buf_1 U13005 ( .ip(n11557), .op(n11617) );
  mux2_1 U13006 ( .ip1(\cache_data[6][3] ), .ip2(n11617), .s(n11496), .op(
        n6060) );
  buf_1 U13007 ( .ip(n11558), .op(n11618) );
  mux2_1 U13008 ( .ip1(\cache_data[6][4] ), .ip2(n11618), .s(n11496), .op(
        n6059) );
  buf_1 U13009 ( .ip(n11559), .op(n11619) );
  mux2_1 U13010 ( .ip1(\cache_data[6][5] ), .ip2(n11619), .s(n11496), .op(
        n6058) );
  buf_1 U13011 ( .ip(n11560), .op(n11620) );
  mux2_1 U13012 ( .ip1(\cache_data[6][6] ), .ip2(n11620), .s(n11496), .op(
        n6057) );
  buf_1 U13013 ( .ip(n11561), .op(n11621) );
  mux2_1 U13014 ( .ip1(\cache_data[6][7] ), .ip2(n11621), .s(n11496), .op(
        n6056) );
  buf_1 U13015 ( .ip(n11562), .op(n11622) );
  mux2_1 U13016 ( .ip1(\cache_data[6][8] ), .ip2(n11622), .s(n11496), .op(
        n6055) );
  buf_1 U13017 ( .ip(n11563), .op(n11623) );
  mux2_1 U13018 ( .ip1(\cache_data[6][9] ), .ip2(n11623), .s(n11496), .op(
        n6054) );
  buf_1 U13019 ( .ip(n11564), .op(n11624) );
  mux2_1 U13020 ( .ip1(\cache_data[6][10] ), .ip2(n11624), .s(n11496), .op(
        n6053) );
  buf_1 U13021 ( .ip(n11565), .op(n11625) );
  mux2_1 U13022 ( .ip1(\cache_data[6][11] ), .ip2(n11625), .s(n11496), .op(
        n6052) );
  buf_1 U13023 ( .ip(n11566), .op(n11626) );
  mux2_1 U13024 ( .ip1(\cache_data[6][12] ), .ip2(n11626), .s(n11496), .op(
        n6051) );
  buf_1 U13025 ( .ip(n11567), .op(n11627) );
  mux2_1 U13026 ( .ip1(\cache_data[6][13] ), .ip2(n11627), .s(n11496), .op(
        n6050) );
  buf_1 U13027 ( .ip(n11568), .op(n11628) );
  mux2_1 U13028 ( .ip1(\cache_data[6][14] ), .ip2(n11628), .s(n11496), .op(
        n6049) );
  buf_1 U13029 ( .ip(n11569), .op(n11629) );
  mux2_1 U13030 ( .ip1(\cache_data[6][15] ), .ip2(n11629), .s(n11496), .op(
        n6048) );
  buf_1 U13031 ( .ip(n11570), .op(n11630) );
  mux2_1 U13032 ( .ip1(\cache_data[6][16] ), .ip2(n11630), .s(n11496), .op(
        n6047) );
  buf_1 U13033 ( .ip(n11571), .op(n11631) );
  mux2_1 U13034 ( .ip1(\cache_data[6][17] ), .ip2(n11631), .s(n11496), .op(
        n6046) );
  buf_1 U13035 ( .ip(n11572), .op(n11632) );
  mux2_1 U13036 ( .ip1(\cache_data[6][18] ), .ip2(n11632), .s(n11496), .op(
        n6045) );
  buf_1 U13037 ( .ip(n11573), .op(n11633) );
  buf_1 U13038 ( .ip(n11496), .op(n11497) );
  mux2_1 U13039 ( .ip1(\cache_data[6][19] ), .ip2(n11633), .s(n11497), .op(
        n6044) );
  buf_1 U13040 ( .ip(n11574), .op(n11634) );
  mux2_1 U13041 ( .ip1(\cache_data[6][20] ), .ip2(n11634), .s(n11497), .op(
        n6043) );
  buf_1 U13042 ( .ip(n11575), .op(n11635) );
  mux2_1 U13043 ( .ip1(\cache_data[6][21] ), .ip2(n11635), .s(n11497), .op(
        n6042) );
  buf_1 U13044 ( .ip(n11576), .op(n11636) );
  mux2_1 U13045 ( .ip1(\cache_data[6][22] ), .ip2(n11636), .s(n11497), .op(
        n6041) );
  buf_1 U13046 ( .ip(n11577), .op(n11637) );
  mux2_1 U13047 ( .ip1(\cache_data[6][23] ), .ip2(n11637), .s(n11497), .op(
        n6040) );
  buf_1 U13048 ( .ip(n11578), .op(n11638) );
  mux2_1 U13049 ( .ip1(\cache_data[6][24] ), .ip2(n11638), .s(n11496), .op(
        n6039) );
  buf_1 U13050 ( .ip(n11580), .op(n11640) );
  mux2_1 U13051 ( .ip1(\cache_data[6][25] ), .ip2(n11640), .s(n11496), .op(
        n6038) );
  buf_1 U13052 ( .ip(n11581), .op(n11641) );
  mux2_1 U13053 ( .ip1(\cache_data[6][26] ), .ip2(n11641), .s(n11497), .op(
        n6037) );
  buf_1 U13054 ( .ip(n11582), .op(n11642) );
  mux2_1 U13055 ( .ip1(\cache_data[6][27] ), .ip2(n11642), .s(n11497), .op(
        n6036) );
  buf_1 U13056 ( .ip(n11583), .op(n11643) );
  mux2_1 U13057 ( .ip1(\cache_data[6][28] ), .ip2(n11643), .s(n11497), .op(
        n6035) );
  buf_1 U13058 ( .ip(n11584), .op(n11644) );
  mux2_1 U13059 ( .ip1(\cache_data[6][29] ), .ip2(n11644), .s(n11497), .op(
        n6034) );
  buf_1 U13060 ( .ip(n11585), .op(n11645) );
  mux2_1 U13061 ( .ip1(\cache_data[6][30] ), .ip2(n11645), .s(n11497), .op(
        n6033) );
  buf_1 U13062 ( .ip(n11587), .op(n11647) );
  mux2_1 U13063 ( .ip1(\cache_data[6][31] ), .ip2(n11647), .s(n11497), .op(
        n6032) );
  nor2_1 U13064 ( .ip1(n11606), .ip2(n11502), .op(n11498) );
  mux2_1 U13065 ( .ip1(\cache_data[6][32] ), .ip2(n11614), .s(n11498), .op(
        n6031) );
  mux2_1 U13066 ( .ip1(\cache_data[6][33] ), .ip2(n11615), .s(n11498), .op(
        n6030) );
  mux2_1 U13067 ( .ip1(\cache_data[6][34] ), .ip2(n11616), .s(n11498), .op(
        n6029) );
  mux2_1 U13068 ( .ip1(\cache_data[6][35] ), .ip2(n11617), .s(n11498), .op(
        n6028) );
  mux2_1 U13069 ( .ip1(\cache_data[6][36] ), .ip2(n11618), .s(n11498), .op(
        n6027) );
  mux2_1 U13070 ( .ip1(\cache_data[6][37] ), .ip2(n11619), .s(n11498), .op(
        n6026) );
  mux2_1 U13071 ( .ip1(\cache_data[6][38] ), .ip2(n11620), .s(n11498), .op(
        n6025) );
  mux2_1 U13072 ( .ip1(\cache_data[6][39] ), .ip2(n11621), .s(n11498), .op(
        n6024) );
  mux2_1 U13073 ( .ip1(\cache_data[6][40] ), .ip2(n11622), .s(n11498), .op(
        n6023) );
  mux2_1 U13074 ( .ip1(\cache_data[6][41] ), .ip2(n11623), .s(n11498), .op(
        n6022) );
  mux2_1 U13075 ( .ip1(\cache_data[6][42] ), .ip2(n11624), .s(n11498), .op(
        n6021) );
  mux2_1 U13076 ( .ip1(\cache_data[6][43] ), .ip2(n11625), .s(n11498), .op(
        n6020) );
  mux2_1 U13077 ( .ip1(\cache_data[6][44] ), .ip2(n11626), .s(n11498), .op(
        n6019) );
  mux2_1 U13078 ( .ip1(\cache_data[6][45] ), .ip2(n11627), .s(n11498), .op(
        n6018) );
  mux2_1 U13079 ( .ip1(\cache_data[6][46] ), .ip2(n11628), .s(n11498), .op(
        n6017) );
  mux2_1 U13080 ( .ip1(\cache_data[6][47] ), .ip2(n11629), .s(n11498), .op(
        n6016) );
  mux2_1 U13081 ( .ip1(\cache_data[6][48] ), .ip2(n11630), .s(n11498), .op(
        n6015) );
  mux2_1 U13082 ( .ip1(\cache_data[6][49] ), .ip2(n11631), .s(n11498), .op(
        n6014) );
  mux2_1 U13083 ( .ip1(\cache_data[6][50] ), .ip2(n11632), .s(n11498), .op(
        n6013) );
  buf_1 U13084 ( .ip(n11498), .op(n11499) );
  mux2_1 U13085 ( .ip1(\cache_data[6][51] ), .ip2(n11633), .s(n11499), .op(
        n6012) );
  mux2_1 U13086 ( .ip1(\cache_data[6][52] ), .ip2(n11634), .s(n11499), .op(
        n6011) );
  mux2_1 U13087 ( .ip1(\cache_data[6][53] ), .ip2(n11635), .s(n11499), .op(
        n6010) );
  mux2_1 U13088 ( .ip1(\cache_data[6][54] ), .ip2(n11636), .s(n11499), .op(
        n6009) );
  mux2_1 U13089 ( .ip1(\cache_data[6][55] ), .ip2(n11637), .s(n11499), .op(
        n6008) );
  mux2_1 U13090 ( .ip1(\cache_data[6][56] ), .ip2(n11638), .s(n11498), .op(
        n6007) );
  mux2_1 U13091 ( .ip1(\cache_data[6][57] ), .ip2(n11640), .s(n11498), .op(
        n6006) );
  mux2_1 U13092 ( .ip1(\cache_data[6][58] ), .ip2(n11641), .s(n11499), .op(
        n6005) );
  mux2_1 U13093 ( .ip1(\cache_data[6][59] ), .ip2(n11642), .s(n11499), .op(
        n6004) );
  mux2_1 U13094 ( .ip1(\cache_data[6][60] ), .ip2(n11643), .s(n11499), .op(
        n6003) );
  mux2_1 U13095 ( .ip1(\cache_data[6][61] ), .ip2(n11644), .s(n11499), .op(
        n6002) );
  mux2_1 U13096 ( .ip1(\cache_data[6][62] ), .ip2(n11645), .s(n11499), .op(
        n6001) );
  mux2_1 U13097 ( .ip1(\cache_data[6][63] ), .ip2(n11647), .s(n11499), .op(
        n6000) );
  nor2_1 U13098 ( .ip1(n11609), .ip2(n11502), .op(n11500) );
  mux2_1 U13099 ( .ip1(\cache_data[6][64] ), .ip2(n11614), .s(n11500), .op(
        n5999) );
  mux2_1 U13100 ( .ip1(\cache_data[6][65] ), .ip2(n11615), .s(n11500), .op(
        n5998) );
  mux2_1 U13101 ( .ip1(\cache_data[6][66] ), .ip2(n11616), .s(n11500), .op(
        n5997) );
  mux2_1 U13102 ( .ip1(\cache_data[6][67] ), .ip2(n11617), .s(n11500), .op(
        n5996) );
  mux2_1 U13103 ( .ip1(\cache_data[6][68] ), .ip2(n11618), .s(n11500), .op(
        n5995) );
  mux2_1 U13104 ( .ip1(\cache_data[6][69] ), .ip2(n11619), .s(n11500), .op(
        n5994) );
  mux2_1 U13105 ( .ip1(\cache_data[6][70] ), .ip2(n11620), .s(n11500), .op(
        n5993) );
  mux2_1 U13106 ( .ip1(\cache_data[6][71] ), .ip2(n11621), .s(n11500), .op(
        n5992) );
  mux2_1 U13107 ( .ip1(\cache_data[6][72] ), .ip2(n11622), .s(n11500), .op(
        n5991) );
  mux2_1 U13108 ( .ip1(\cache_data[6][73] ), .ip2(n11623), .s(n11500), .op(
        n5990) );
  mux2_1 U13109 ( .ip1(\cache_data[6][74] ), .ip2(n11624), .s(n11500), .op(
        n5989) );
  mux2_1 U13110 ( .ip1(\cache_data[6][75] ), .ip2(n11625), .s(n11500), .op(
        n5988) );
  mux2_1 U13111 ( .ip1(\cache_data[6][76] ), .ip2(n11626), .s(n11500), .op(
        n5987) );
  mux2_1 U13112 ( .ip1(\cache_data[6][77] ), .ip2(n11627), .s(n11500), .op(
        n5986) );
  mux2_1 U13113 ( .ip1(\cache_data[6][78] ), .ip2(n11628), .s(n11500), .op(
        n5985) );
  mux2_1 U13114 ( .ip1(\cache_data[6][79] ), .ip2(n11629), .s(n11500), .op(
        n5984) );
  mux2_1 U13115 ( .ip1(\cache_data[6][80] ), .ip2(n11630), .s(n11500), .op(
        n5983) );
  mux2_1 U13116 ( .ip1(\cache_data[6][81] ), .ip2(n11631), .s(n11500), .op(
        n5982) );
  mux2_1 U13117 ( .ip1(\cache_data[6][82] ), .ip2(n11632), .s(n11500), .op(
        n5981) );
  buf_1 U13118 ( .ip(n11500), .op(n11501) );
  mux2_1 U13119 ( .ip1(\cache_data[6][83] ), .ip2(n11633), .s(n11501), .op(
        n5980) );
  mux2_1 U13120 ( .ip1(\cache_data[6][84] ), .ip2(n11634), .s(n11501), .op(
        n5979) );
  mux2_1 U13121 ( .ip1(\cache_data[6][85] ), .ip2(n11635), .s(n11501), .op(
        n5978) );
  mux2_1 U13122 ( .ip1(\cache_data[6][86] ), .ip2(n11636), .s(n11501), .op(
        n5977) );
  mux2_1 U13123 ( .ip1(\cache_data[6][87] ), .ip2(n11637), .s(n11501), .op(
        n5976) );
  mux2_1 U13124 ( .ip1(\cache_data[6][88] ), .ip2(n11638), .s(n11500), .op(
        n5975) );
  mux2_1 U13125 ( .ip1(\cache_data[6][89] ), .ip2(n11640), .s(n11500), .op(
        n5974) );
  mux2_1 U13126 ( .ip1(\cache_data[6][90] ), .ip2(n11641), .s(n11501), .op(
        n5973) );
  mux2_1 U13127 ( .ip1(\cache_data[6][91] ), .ip2(n11642), .s(n11501), .op(
        n5972) );
  mux2_1 U13128 ( .ip1(\cache_data[6][92] ), .ip2(n11643), .s(n11501), .op(
        n5971) );
  mux2_1 U13129 ( .ip1(\cache_data[6][93] ), .ip2(n11644), .s(n11501), .op(
        n5970) );
  mux2_1 U13130 ( .ip1(\cache_data[6][94] ), .ip2(n11645), .s(n11501), .op(
        n5969) );
  mux2_1 U13131 ( .ip1(\cache_data[6][95] ), .ip2(n11647), .s(n11501), .op(
        n5968) );
  nor2_1 U13132 ( .ip1(n11613), .ip2(n11502), .op(n11503) );
  mux2_1 U13133 ( .ip1(\cache_data[6][96] ), .ip2(n11614), .s(n11503), .op(
        n5967) );
  mux2_1 U13134 ( .ip1(\cache_data[6][97] ), .ip2(n11615), .s(n11503), .op(
        n5966) );
  mux2_1 U13135 ( .ip1(\cache_data[6][98] ), .ip2(n11616), .s(n11503), .op(
        n5965) );
  mux2_1 U13136 ( .ip1(\cache_data[6][99] ), .ip2(n11617), .s(n11503), .op(
        n5964) );
  mux2_1 U13137 ( .ip1(\cache_data[6][100] ), .ip2(n11618), .s(n11503), .op(
        n5963) );
  mux2_1 U13138 ( .ip1(\cache_data[6][101] ), .ip2(n11619), .s(n11503), .op(
        n5962) );
  mux2_1 U13139 ( .ip1(\cache_data[6][102] ), .ip2(n11620), .s(n11503), .op(
        n5961) );
  mux2_1 U13140 ( .ip1(\cache_data[6][103] ), .ip2(n11621), .s(n11503), .op(
        n5960) );
  mux2_1 U13141 ( .ip1(\cache_data[6][104] ), .ip2(n11622), .s(n11503), .op(
        n5959) );
  mux2_1 U13142 ( .ip1(\cache_data[6][105] ), .ip2(n11623), .s(n11503), .op(
        n5958) );
  mux2_1 U13143 ( .ip1(\cache_data[6][106] ), .ip2(n11624), .s(n11503), .op(
        n5957) );
  mux2_1 U13144 ( .ip1(\cache_data[6][107] ), .ip2(n11625), .s(n11503), .op(
        n5956) );
  mux2_1 U13145 ( .ip1(\cache_data[6][108] ), .ip2(n11626), .s(n11503), .op(
        n5955) );
  mux2_1 U13146 ( .ip1(\cache_data[6][109] ), .ip2(n11627), .s(n11503), .op(
        n5954) );
  mux2_1 U13147 ( .ip1(\cache_data[6][110] ), .ip2(n11628), .s(n11503), .op(
        n5953) );
  mux2_1 U13148 ( .ip1(\cache_data[6][111] ), .ip2(n11629), .s(n11503), .op(
        n5952) );
  mux2_1 U13149 ( .ip1(\cache_data[6][112] ), .ip2(n11630), .s(n11503), .op(
        n5951) );
  mux2_1 U13150 ( .ip1(\cache_data[6][113] ), .ip2(n11631), .s(n11503), .op(
        n5950) );
  mux2_1 U13151 ( .ip1(\cache_data[6][114] ), .ip2(n11632), .s(n11503), .op(
        n5949) );
  buf_1 U13152 ( .ip(n11503), .op(n11504) );
  mux2_1 U13153 ( .ip1(\cache_data[6][115] ), .ip2(n11633), .s(n11504), .op(
        n5948) );
  mux2_1 U13154 ( .ip1(\cache_data[6][116] ), .ip2(n11634), .s(n11504), .op(
        n5947) );
  mux2_1 U13155 ( .ip1(\cache_data[6][117] ), .ip2(n11635), .s(n11504), .op(
        n5946) );
  mux2_1 U13156 ( .ip1(\cache_data[6][118] ), .ip2(n11636), .s(n11504), .op(
        n5945) );
  mux2_1 U13157 ( .ip1(\cache_data[6][119] ), .ip2(n11637), .s(n11504), .op(
        n5944) );
  mux2_1 U13158 ( .ip1(\cache_data[6][120] ), .ip2(n11638), .s(n11503), .op(
        n5943) );
  mux2_1 U13159 ( .ip1(\cache_data[6][121] ), .ip2(n11640), .s(n11503), .op(
        n5942) );
  mux2_1 U13160 ( .ip1(\cache_data[6][122] ), .ip2(n11641), .s(n11504), .op(
        n5941) );
  mux2_1 U13161 ( .ip1(\cache_data[6][123] ), .ip2(n11642), .s(n11504), .op(
        n5940) );
  mux2_1 U13162 ( .ip1(\cache_data[6][124] ), .ip2(n11643), .s(n11504), .op(
        n5939) );
  mux2_1 U13163 ( .ip1(\cache_data[6][125] ), .ip2(n11644), .s(n11504), .op(
        n5938) );
  mux2_1 U13164 ( .ip1(\cache_data[6][126] ), .ip2(n11645), .s(n11504), .op(
        n5937) );
  mux2_1 U13165 ( .ip1(\cache_data[6][127] ), .ip2(n11647), .s(n11504), .op(
        n5936) );
  nor2_1 U13166 ( .ip1(n11603), .ip2(n8153), .op(n11505) );
  mux2_1 U13167 ( .ip1(\cache_data[7][0] ), .ip2(n11614), .s(n11505), .op(
        n5935) );
  mux2_1 U13168 ( .ip1(\cache_data[7][1] ), .ip2(n11615), .s(n11505), .op(
        n5934) );
  mux2_1 U13169 ( .ip1(\cache_data[7][2] ), .ip2(n11616), .s(n11505), .op(
        n5933) );
  mux2_1 U13170 ( .ip1(\cache_data[7][3] ), .ip2(n11617), .s(n11505), .op(
        n5932) );
  mux2_1 U13171 ( .ip1(\cache_data[7][4] ), .ip2(n11618), .s(n11505), .op(
        n5931) );
  mux2_1 U13172 ( .ip1(\cache_data[7][5] ), .ip2(n11619), .s(n11505), .op(
        n5930) );
  mux2_1 U13173 ( .ip1(\cache_data[7][6] ), .ip2(n11620), .s(n11505), .op(
        n5929) );
  mux2_1 U13174 ( .ip1(\cache_data[7][7] ), .ip2(n11621), .s(n11505), .op(
        n5928) );
  mux2_1 U13175 ( .ip1(\cache_data[7][8] ), .ip2(n11622), .s(n11505), .op(
        n5927) );
  mux2_1 U13176 ( .ip1(\cache_data[7][9] ), .ip2(n11623), .s(n11505), .op(
        n5926) );
  mux2_1 U13177 ( .ip1(\cache_data[7][10] ), .ip2(n11624), .s(n11505), .op(
        n5925) );
  mux2_1 U13178 ( .ip1(\cache_data[7][11] ), .ip2(n11625), .s(n11505), .op(
        n5924) );
  mux2_1 U13179 ( .ip1(\cache_data[7][12] ), .ip2(n11626), .s(n11505), .op(
        n5923) );
  mux2_1 U13180 ( .ip1(\cache_data[7][13] ), .ip2(n11627), .s(n11505), .op(
        n5922) );
  mux2_1 U13181 ( .ip1(\cache_data[7][14] ), .ip2(n11628), .s(n11505), .op(
        n5921) );
  mux2_1 U13182 ( .ip1(\cache_data[7][15] ), .ip2(n11629), .s(n11505), .op(
        n5920) );
  mux2_1 U13183 ( .ip1(\cache_data[7][16] ), .ip2(n11630), .s(n11505), .op(
        n5919) );
  mux2_1 U13184 ( .ip1(\cache_data[7][17] ), .ip2(n11631), .s(n11505), .op(
        n5918) );
  mux2_1 U13185 ( .ip1(\cache_data[7][18] ), .ip2(n11632), .s(n11505), .op(
        n5917) );
  buf_1 U13186 ( .ip(n11505), .op(n11506) );
  mux2_1 U13187 ( .ip1(\cache_data[7][19] ), .ip2(n11633), .s(n11506), .op(
        n5916) );
  mux2_1 U13188 ( .ip1(\cache_data[7][20] ), .ip2(n11634), .s(n11506), .op(
        n5915) );
  mux2_1 U13189 ( .ip1(\cache_data[7][21] ), .ip2(n11635), .s(n11506), .op(
        n5914) );
  mux2_1 U13190 ( .ip1(\cache_data[7][22] ), .ip2(n11636), .s(n11506), .op(
        n5913) );
  mux2_1 U13191 ( .ip1(\cache_data[7][23] ), .ip2(n11637), .s(n11506), .op(
        n5912) );
  mux2_1 U13192 ( .ip1(\cache_data[7][24] ), .ip2(n11638), .s(n11505), .op(
        n5911) );
  mux2_1 U13193 ( .ip1(\cache_data[7][25] ), .ip2(n11640), .s(n11505), .op(
        n5910) );
  mux2_1 U13194 ( .ip1(\cache_data[7][26] ), .ip2(n11641), .s(n11506), .op(
        n5909) );
  mux2_1 U13195 ( .ip1(\cache_data[7][27] ), .ip2(n11642), .s(n11506), .op(
        n5908) );
  mux2_1 U13196 ( .ip1(\cache_data[7][28] ), .ip2(n11643), .s(n11506), .op(
        n5907) );
  mux2_1 U13197 ( .ip1(\cache_data[7][29] ), .ip2(n11644), .s(n11506), .op(
        n5906) );
  mux2_1 U13198 ( .ip1(\cache_data[7][30] ), .ip2(n11645), .s(n11506), .op(
        n5905) );
  mux2_1 U13199 ( .ip1(\cache_data[7][31] ), .ip2(n11647), .s(n11506), .op(
        n5904) );
  nor2_1 U13200 ( .ip1(n11606), .ip2(n8153), .op(n11507) );
  mux2_1 U13201 ( .ip1(\cache_data[7][32] ), .ip2(n11614), .s(n11507), .op(
        n5903) );
  mux2_1 U13202 ( .ip1(\cache_data[7][33] ), .ip2(n11615), .s(n11507), .op(
        n5902) );
  mux2_1 U13203 ( .ip1(\cache_data[7][34] ), .ip2(n11616), .s(n11507), .op(
        n5901) );
  mux2_1 U13204 ( .ip1(\cache_data[7][35] ), .ip2(n11617), .s(n11507), .op(
        n5900) );
  mux2_1 U13205 ( .ip1(\cache_data[7][36] ), .ip2(n11618), .s(n11507), .op(
        n5899) );
  mux2_1 U13206 ( .ip1(\cache_data[7][37] ), .ip2(n11619), .s(n11507), .op(
        n5898) );
  mux2_1 U13207 ( .ip1(\cache_data[7][38] ), .ip2(n11620), .s(n11507), .op(
        n5897) );
  mux2_1 U13208 ( .ip1(\cache_data[7][39] ), .ip2(n11621), .s(n11507), .op(
        n5896) );
  mux2_1 U13209 ( .ip1(\cache_data[7][40] ), .ip2(n11622), .s(n11507), .op(
        n5895) );
  mux2_1 U13210 ( .ip1(\cache_data[7][41] ), .ip2(n11623), .s(n11507), .op(
        n5894) );
  mux2_1 U13211 ( .ip1(\cache_data[7][42] ), .ip2(n11624), .s(n11507), .op(
        n5893) );
  mux2_1 U13212 ( .ip1(\cache_data[7][43] ), .ip2(n11625), .s(n11507), .op(
        n5892) );
  mux2_1 U13213 ( .ip1(\cache_data[7][44] ), .ip2(n11626), .s(n11507), .op(
        n5891) );
  mux2_1 U13214 ( .ip1(\cache_data[7][45] ), .ip2(n11627), .s(n11507), .op(
        n5890) );
  mux2_1 U13215 ( .ip1(\cache_data[7][46] ), .ip2(n11628), .s(n11507), .op(
        n5889) );
  mux2_1 U13216 ( .ip1(\cache_data[7][47] ), .ip2(n11629), .s(n11507), .op(
        n5888) );
  mux2_1 U13217 ( .ip1(\cache_data[7][48] ), .ip2(n11630), .s(n11507), .op(
        n5887) );
  mux2_1 U13218 ( .ip1(\cache_data[7][49] ), .ip2(n11631), .s(n11507), .op(
        n5886) );
  mux2_1 U13219 ( .ip1(\cache_data[7][50] ), .ip2(n11632), .s(n11507), .op(
        n5885) );
  buf_1 U13220 ( .ip(n11507), .op(n11508) );
  mux2_1 U13221 ( .ip1(\cache_data[7][51] ), .ip2(n11633), .s(n11508), .op(
        n5884) );
  mux2_1 U13222 ( .ip1(\cache_data[7][52] ), .ip2(n11634), .s(n11508), .op(
        n5883) );
  mux2_1 U13223 ( .ip1(\cache_data[7][53] ), .ip2(n11635), .s(n11508), .op(
        n5882) );
  mux2_1 U13224 ( .ip1(\cache_data[7][54] ), .ip2(n11636), .s(n11508), .op(
        n5881) );
  mux2_1 U13225 ( .ip1(\cache_data[7][55] ), .ip2(n11637), .s(n11508), .op(
        n5880) );
  mux2_1 U13226 ( .ip1(\cache_data[7][56] ), .ip2(n11638), .s(n11507), .op(
        n5879) );
  mux2_1 U13227 ( .ip1(\cache_data[7][57] ), .ip2(n11640), .s(n11507), .op(
        n5878) );
  mux2_1 U13228 ( .ip1(\cache_data[7][58] ), .ip2(n11641), .s(n11508), .op(
        n5877) );
  mux2_1 U13229 ( .ip1(\cache_data[7][59] ), .ip2(n11642), .s(n11508), .op(
        n5876) );
  mux2_1 U13230 ( .ip1(\cache_data[7][60] ), .ip2(n11643), .s(n11508), .op(
        n5875) );
  mux2_1 U13231 ( .ip1(\cache_data[7][61] ), .ip2(n11644), .s(n11508), .op(
        n5874) );
  mux2_1 U13232 ( .ip1(\cache_data[7][62] ), .ip2(n11645), .s(n11508), .op(
        n5873) );
  mux2_1 U13233 ( .ip1(\cache_data[7][63] ), .ip2(n11647), .s(n11508), .op(
        n5872) );
  nor2_1 U13234 ( .ip1(n11609), .ip2(n8153), .op(n11509) );
  mux2_1 U13235 ( .ip1(\cache_data[7][64] ), .ip2(n11614), .s(n11509), .op(
        n5871) );
  mux2_1 U13236 ( .ip1(\cache_data[7][65] ), .ip2(n11615), .s(n11509), .op(
        n5870) );
  mux2_1 U13237 ( .ip1(\cache_data[7][66] ), .ip2(n11616), .s(n11509), .op(
        n5869) );
  mux2_1 U13238 ( .ip1(\cache_data[7][67] ), .ip2(n11617), .s(n11509), .op(
        n5868) );
  mux2_1 U13239 ( .ip1(\cache_data[7][68] ), .ip2(n11618), .s(n11509), .op(
        n5867) );
  mux2_1 U13240 ( .ip1(\cache_data[7][69] ), .ip2(n11619), .s(n11509), .op(
        n5866) );
  mux2_1 U13241 ( .ip1(\cache_data[7][70] ), .ip2(n11620), .s(n11509), .op(
        n5865) );
  mux2_1 U13242 ( .ip1(\cache_data[7][71] ), .ip2(n11621), .s(n11509), .op(
        n5864) );
  mux2_1 U13243 ( .ip1(\cache_data[7][72] ), .ip2(n11622), .s(n11509), .op(
        n5863) );
  mux2_1 U13244 ( .ip1(\cache_data[7][73] ), .ip2(n11623), .s(n11509), .op(
        n5862) );
  mux2_1 U13245 ( .ip1(\cache_data[7][74] ), .ip2(n11624), .s(n11509), .op(
        n5861) );
  mux2_1 U13246 ( .ip1(\cache_data[7][75] ), .ip2(n11625), .s(n11509), .op(
        n5860) );
  mux2_1 U13247 ( .ip1(\cache_data[7][76] ), .ip2(n11626), .s(n11509), .op(
        n5859) );
  mux2_1 U13248 ( .ip1(\cache_data[7][77] ), .ip2(n11627), .s(n11509), .op(
        n5858) );
  mux2_1 U13249 ( .ip1(\cache_data[7][78] ), .ip2(n11628), .s(n11509), .op(
        n5857) );
  mux2_1 U13250 ( .ip1(\cache_data[7][79] ), .ip2(n11629), .s(n11509), .op(
        n5856) );
  mux2_1 U13251 ( .ip1(\cache_data[7][80] ), .ip2(n11630), .s(n11509), .op(
        n5855) );
  mux2_1 U13252 ( .ip1(\cache_data[7][81] ), .ip2(n11631), .s(n11509), .op(
        n5854) );
  mux2_1 U13253 ( .ip1(\cache_data[7][82] ), .ip2(n11632), .s(n11509), .op(
        n5853) );
  buf_1 U13254 ( .ip(n11509), .op(n11510) );
  mux2_1 U13255 ( .ip1(\cache_data[7][83] ), .ip2(n11633), .s(n11510), .op(
        n5852) );
  mux2_1 U13256 ( .ip1(\cache_data[7][84] ), .ip2(n11634), .s(n11510), .op(
        n5851) );
  mux2_1 U13257 ( .ip1(\cache_data[7][85] ), .ip2(n11635), .s(n11510), .op(
        n5850) );
  mux2_1 U13258 ( .ip1(\cache_data[7][86] ), .ip2(n11636), .s(n11510), .op(
        n5849) );
  mux2_1 U13259 ( .ip1(\cache_data[7][87] ), .ip2(n11637), .s(n11510), .op(
        n5848) );
  mux2_1 U13260 ( .ip1(\cache_data[7][88] ), .ip2(n11638), .s(n11509), .op(
        n5847) );
  mux2_1 U13261 ( .ip1(\cache_data[7][89] ), .ip2(n11640), .s(n11509), .op(
        n5846) );
  mux2_1 U13262 ( .ip1(\cache_data[7][90] ), .ip2(n11641), .s(n11510), .op(
        n5845) );
  mux2_1 U13263 ( .ip1(\cache_data[7][91] ), .ip2(n11642), .s(n11510), .op(
        n5844) );
  mux2_1 U13264 ( .ip1(\cache_data[7][92] ), .ip2(n11643), .s(n11510), .op(
        n5843) );
  mux2_1 U13265 ( .ip1(\cache_data[7][93] ), .ip2(n11644), .s(n11510), .op(
        n5842) );
  mux2_1 U13266 ( .ip1(\cache_data[7][94] ), .ip2(n11645), .s(n11510), .op(
        n5841) );
  mux2_1 U13267 ( .ip1(\cache_data[7][95] ), .ip2(n11647), .s(n11510), .op(
        n5840) );
  nor2_1 U13268 ( .ip1(n11613), .ip2(n8153), .op(n11511) );
  mux2_1 U13269 ( .ip1(\cache_data[7][96] ), .ip2(n11614), .s(n11511), .op(
        n5839) );
  mux2_1 U13270 ( .ip1(\cache_data[7][97] ), .ip2(n11615), .s(n11511), .op(
        n5838) );
  mux2_1 U13271 ( .ip1(\cache_data[7][98] ), .ip2(n11616), .s(n11511), .op(
        n5837) );
  mux2_1 U13272 ( .ip1(\cache_data[7][99] ), .ip2(n11617), .s(n11511), .op(
        n5836) );
  mux2_1 U13273 ( .ip1(\cache_data[7][100] ), .ip2(n11618), .s(n11511), .op(
        n5835) );
  mux2_1 U13274 ( .ip1(\cache_data[7][101] ), .ip2(n11619), .s(n11511), .op(
        n5834) );
  mux2_1 U13275 ( .ip1(\cache_data[7][102] ), .ip2(n11620), .s(n11511), .op(
        n5833) );
  mux2_1 U13276 ( .ip1(\cache_data[7][103] ), .ip2(n11621), .s(n11511), .op(
        n5832) );
  mux2_1 U13277 ( .ip1(\cache_data[7][104] ), .ip2(n11622), .s(n11511), .op(
        n5831) );
  mux2_1 U13278 ( .ip1(\cache_data[7][105] ), .ip2(n11623), .s(n11511), .op(
        n5830) );
  mux2_1 U13279 ( .ip1(\cache_data[7][106] ), .ip2(n11624), .s(n11511), .op(
        n5829) );
  mux2_1 U13280 ( .ip1(\cache_data[7][107] ), .ip2(n11625), .s(n11511), .op(
        n5828) );
  mux2_1 U13281 ( .ip1(\cache_data[7][108] ), .ip2(n11626), .s(n11511), .op(
        n5827) );
  mux2_1 U13282 ( .ip1(\cache_data[7][109] ), .ip2(n11627), .s(n11511), .op(
        n5826) );
  mux2_1 U13283 ( .ip1(\cache_data[7][110] ), .ip2(n11628), .s(n11511), .op(
        n5825) );
  mux2_1 U13284 ( .ip1(\cache_data[7][111] ), .ip2(n11629), .s(n11511), .op(
        n5824) );
  mux2_1 U13285 ( .ip1(\cache_data[7][112] ), .ip2(n11630), .s(n11511), .op(
        n5823) );
  mux2_1 U13286 ( .ip1(\cache_data[7][113] ), .ip2(n11631), .s(n11511), .op(
        n5822) );
  mux2_1 U13287 ( .ip1(\cache_data[7][114] ), .ip2(n11632), .s(n11511), .op(
        n5821) );
  buf_1 U13288 ( .ip(n11511), .op(n11512) );
  mux2_1 U13289 ( .ip1(\cache_data[7][115] ), .ip2(n11633), .s(n11512), .op(
        n5820) );
  mux2_1 U13290 ( .ip1(\cache_data[7][116] ), .ip2(n11634), .s(n11512), .op(
        n5819) );
  mux2_1 U13291 ( .ip1(\cache_data[7][117] ), .ip2(n11635), .s(n11512), .op(
        n5818) );
  mux2_1 U13292 ( .ip1(\cache_data[7][118] ), .ip2(n11636), .s(n11512), .op(
        n5817) );
  mux2_1 U13293 ( .ip1(\cache_data[7][119] ), .ip2(n11637), .s(n11512), .op(
        n5816) );
  mux2_1 U13294 ( .ip1(\cache_data[7][120] ), .ip2(n11638), .s(n11511), .op(
        n5815) );
  mux2_1 U13295 ( .ip1(\cache_data[7][121] ), .ip2(n11640), .s(n11511), .op(
        n5814) );
  mux2_1 U13296 ( .ip1(\cache_data[7][122] ), .ip2(n11641), .s(n11512), .op(
        n5813) );
  mux2_1 U13297 ( .ip1(\cache_data[7][123] ), .ip2(n11642), .s(n11512), .op(
        n5812) );
  mux2_1 U13298 ( .ip1(\cache_data[7][124] ), .ip2(n11643), .s(n11512), .op(
        n5811) );
  mux2_1 U13299 ( .ip1(\cache_data[7][125] ), .ip2(n11644), .s(n11512), .op(
        n5810) );
  mux2_1 U13300 ( .ip1(\cache_data[7][126] ), .ip2(n11645), .s(n11512), .op(
        n5809) );
  mux2_1 U13301 ( .ip1(\cache_data[7][127] ), .ip2(n11647), .s(n11512), .op(
        n5808) );
  nor2_1 U13302 ( .ip1(n11603), .ip2(n8137), .op(n11513) );
  mux2_1 U13303 ( .ip1(\cache_data[8][0] ), .ip2(n11554), .s(n11513), .op(
        n5807) );
  mux2_1 U13304 ( .ip1(\cache_data[8][1] ), .ip2(n11555), .s(n11513), .op(
        n5806) );
  mux2_1 U13305 ( .ip1(\cache_data[8][2] ), .ip2(n11556), .s(n11513), .op(
        n5805) );
  mux2_1 U13306 ( .ip1(\cache_data[8][3] ), .ip2(n11557), .s(n11513), .op(
        n5804) );
  mux2_1 U13307 ( .ip1(\cache_data[8][4] ), .ip2(n11558), .s(n11513), .op(
        n5803) );
  mux2_1 U13308 ( .ip1(\cache_data[8][5] ), .ip2(n11559), .s(n11513), .op(
        n5802) );
  mux2_1 U13309 ( .ip1(\cache_data[8][6] ), .ip2(n11560), .s(n11513), .op(
        n5801) );
  mux2_1 U13310 ( .ip1(\cache_data[8][7] ), .ip2(n11561), .s(n11513), .op(
        n5800) );
  mux2_1 U13311 ( .ip1(\cache_data[8][8] ), .ip2(n11562), .s(n11513), .op(
        n5799) );
  mux2_1 U13312 ( .ip1(\cache_data[8][9] ), .ip2(n11563), .s(n11513), .op(
        n5798) );
  mux2_1 U13313 ( .ip1(\cache_data[8][10] ), .ip2(n11564), .s(n11513), .op(
        n5797) );
  mux2_1 U13314 ( .ip1(\cache_data[8][11] ), .ip2(n11565), .s(n11513), .op(
        n5796) );
  mux2_1 U13315 ( .ip1(\cache_data[8][12] ), .ip2(n11566), .s(n11513), .op(
        n5795) );
  mux2_1 U13316 ( .ip1(\cache_data[8][13] ), .ip2(n11567), .s(n11513), .op(
        n5794) );
  mux2_1 U13317 ( .ip1(\cache_data[8][14] ), .ip2(n11568), .s(n11513), .op(
        n5793) );
  mux2_1 U13318 ( .ip1(\cache_data[8][15] ), .ip2(n11569), .s(n11513), .op(
        n5792) );
  mux2_1 U13319 ( .ip1(\cache_data[8][16] ), .ip2(n11570), .s(n11513), .op(
        n5791) );
  mux2_1 U13320 ( .ip1(\cache_data[8][17] ), .ip2(n11571), .s(n11513), .op(
        n5790) );
  mux2_1 U13321 ( .ip1(\cache_data[8][18] ), .ip2(n11572), .s(n11513), .op(
        n5789) );
  buf_1 U13322 ( .ip(n11513), .op(n11514) );
  mux2_1 U13323 ( .ip1(\cache_data[8][19] ), .ip2(n11573), .s(n11514), .op(
        n5788) );
  mux2_1 U13324 ( .ip1(\cache_data[8][20] ), .ip2(n11574), .s(n11514), .op(
        n5787) );
  mux2_1 U13325 ( .ip1(\cache_data[8][21] ), .ip2(n11575), .s(n11514), .op(
        n5786) );
  mux2_1 U13326 ( .ip1(\cache_data[8][22] ), .ip2(n11576), .s(n11514), .op(
        n5785) );
  mux2_1 U13327 ( .ip1(\cache_data[8][23] ), .ip2(n11577), .s(n11514), .op(
        n5784) );
  mux2_1 U13328 ( .ip1(\cache_data[8][24] ), .ip2(n11578), .s(n11513), .op(
        n5783) );
  mux2_1 U13329 ( .ip1(\cache_data[8][25] ), .ip2(n11580), .s(n11513), .op(
        n5782) );
  mux2_1 U13330 ( .ip1(\cache_data[8][26] ), .ip2(n11581), .s(n11514), .op(
        n5781) );
  mux2_1 U13331 ( .ip1(\cache_data[8][27] ), .ip2(n11582), .s(n11514), .op(
        n5780) );
  mux2_1 U13332 ( .ip1(\cache_data[8][28] ), .ip2(n11583), .s(n11514), .op(
        n5779) );
  mux2_1 U13333 ( .ip1(\cache_data[8][29] ), .ip2(n11584), .s(n11514), .op(
        n5778) );
  mux2_1 U13334 ( .ip1(\cache_data[8][30] ), .ip2(n11585), .s(n11514), .op(
        n5777) );
  mux2_1 U13335 ( .ip1(\cache_data[8][31] ), .ip2(n11587), .s(n11514), .op(
        n5776) );
  nor2_1 U13336 ( .ip1(n11606), .ip2(n8137), .op(n11515) );
  mux2_1 U13337 ( .ip1(\cache_data[8][32] ), .ip2(n11554), .s(n11515), .op(
        n5775) );
  mux2_1 U13338 ( .ip1(\cache_data[8][33] ), .ip2(n11555), .s(n11515), .op(
        n5774) );
  mux2_1 U13339 ( .ip1(\cache_data[8][34] ), .ip2(n11556), .s(n11515), .op(
        n5773) );
  mux2_1 U13340 ( .ip1(\cache_data[8][35] ), .ip2(n11557), .s(n11515), .op(
        n5772) );
  mux2_1 U13341 ( .ip1(\cache_data[8][36] ), .ip2(n11558), .s(n11515), .op(
        n5771) );
  mux2_1 U13342 ( .ip1(\cache_data[8][37] ), .ip2(n11559), .s(n11515), .op(
        n5770) );
  mux2_1 U13343 ( .ip1(\cache_data[8][38] ), .ip2(n11560), .s(n11515), .op(
        n5769) );
  mux2_1 U13344 ( .ip1(\cache_data[8][39] ), .ip2(n11561), .s(n11515), .op(
        n5768) );
  mux2_1 U13345 ( .ip1(\cache_data[8][40] ), .ip2(n11562), .s(n11515), .op(
        n5767) );
  mux2_1 U13346 ( .ip1(\cache_data[8][41] ), .ip2(n11563), .s(n11515), .op(
        n5766) );
  mux2_1 U13347 ( .ip1(\cache_data[8][42] ), .ip2(n11564), .s(n11515), .op(
        n5765) );
  mux2_1 U13348 ( .ip1(\cache_data[8][43] ), .ip2(n11565), .s(n11515), .op(
        n5764) );
  mux2_1 U13349 ( .ip1(\cache_data[8][44] ), .ip2(n11566), .s(n11515), .op(
        n5763) );
  mux2_1 U13350 ( .ip1(\cache_data[8][45] ), .ip2(n11567), .s(n11515), .op(
        n5762) );
  mux2_1 U13351 ( .ip1(\cache_data[8][46] ), .ip2(n11568), .s(n11515), .op(
        n5761) );
  mux2_1 U13352 ( .ip1(\cache_data[8][47] ), .ip2(n11569), .s(n11515), .op(
        n5760) );
  mux2_1 U13353 ( .ip1(\cache_data[8][48] ), .ip2(n11570), .s(n11515), .op(
        n5759) );
  mux2_1 U13354 ( .ip1(\cache_data[8][49] ), .ip2(n11571), .s(n11515), .op(
        n5758) );
  mux2_1 U13355 ( .ip1(\cache_data[8][50] ), .ip2(n11572), .s(n11515), .op(
        n5757) );
  buf_1 U13356 ( .ip(n11515), .op(n11516) );
  mux2_1 U13357 ( .ip1(\cache_data[8][51] ), .ip2(n11573), .s(n11516), .op(
        n5756) );
  mux2_1 U13358 ( .ip1(\cache_data[8][52] ), .ip2(n11574), .s(n11516), .op(
        n5755) );
  mux2_1 U13359 ( .ip1(\cache_data[8][53] ), .ip2(n11575), .s(n11516), .op(
        n5754) );
  mux2_1 U13360 ( .ip1(\cache_data[8][54] ), .ip2(n11576), .s(n11516), .op(
        n5753) );
  mux2_1 U13361 ( .ip1(\cache_data[8][55] ), .ip2(n11577), .s(n11516), .op(
        n5752) );
  mux2_1 U13362 ( .ip1(\cache_data[8][56] ), .ip2(n11578), .s(n11515), .op(
        n5751) );
  mux2_1 U13363 ( .ip1(\cache_data[8][57] ), .ip2(n11580), .s(n11515), .op(
        n5750) );
  mux2_1 U13364 ( .ip1(\cache_data[8][58] ), .ip2(n11581), .s(n11516), .op(
        n5749) );
  mux2_1 U13365 ( .ip1(\cache_data[8][59] ), .ip2(n11582), .s(n11516), .op(
        n5748) );
  mux2_1 U13366 ( .ip1(\cache_data[8][60] ), .ip2(n11583), .s(n11516), .op(
        n5747) );
  mux2_1 U13367 ( .ip1(\cache_data[8][61] ), .ip2(n11584), .s(n11516), .op(
        n5746) );
  mux2_1 U13368 ( .ip1(\cache_data[8][62] ), .ip2(n11585), .s(n11516), .op(
        n5745) );
  mux2_1 U13369 ( .ip1(\cache_data[8][63] ), .ip2(n11587), .s(n11516), .op(
        n5744) );
  nor2_1 U13370 ( .ip1(n11609), .ip2(n8137), .op(n11517) );
  mux2_1 U13371 ( .ip1(\cache_data[8][64] ), .ip2(n11614), .s(n11517), .op(
        n5743) );
  mux2_1 U13372 ( .ip1(\cache_data[8][65] ), .ip2(n11615), .s(n11517), .op(
        n5742) );
  mux2_1 U13373 ( .ip1(\cache_data[8][66] ), .ip2(n11616), .s(n11517), .op(
        n5741) );
  mux2_1 U13374 ( .ip1(\cache_data[8][67] ), .ip2(n11617), .s(n11517), .op(
        n5740) );
  mux2_1 U13375 ( .ip1(\cache_data[8][68] ), .ip2(n11618), .s(n11517), .op(
        n5739) );
  mux2_1 U13376 ( .ip1(\cache_data[8][69] ), .ip2(n11619), .s(n11517), .op(
        n5738) );
  mux2_1 U13377 ( .ip1(\cache_data[8][70] ), .ip2(n11620), .s(n11517), .op(
        n5737) );
  mux2_1 U13378 ( .ip1(\cache_data[8][71] ), .ip2(n11621), .s(n11517), .op(
        n5736) );
  mux2_1 U13379 ( .ip1(\cache_data[8][72] ), .ip2(n11622), .s(n11517), .op(
        n5735) );
  mux2_1 U13380 ( .ip1(\cache_data[8][73] ), .ip2(n11623), .s(n11517), .op(
        n5734) );
  mux2_1 U13381 ( .ip1(\cache_data[8][74] ), .ip2(n11624), .s(n11517), .op(
        n5733) );
  mux2_1 U13382 ( .ip1(\cache_data[8][75] ), .ip2(n11625), .s(n11517), .op(
        n5732) );
  mux2_1 U13383 ( .ip1(\cache_data[8][76] ), .ip2(n11626), .s(n11517), .op(
        n5731) );
  mux2_1 U13384 ( .ip1(\cache_data[8][77] ), .ip2(n11627), .s(n11517), .op(
        n5730) );
  mux2_1 U13385 ( .ip1(\cache_data[8][78] ), .ip2(n11628), .s(n11517), .op(
        n5729) );
  mux2_1 U13386 ( .ip1(\cache_data[8][79] ), .ip2(n11629), .s(n11517), .op(
        n5728) );
  mux2_1 U13387 ( .ip1(\cache_data[8][80] ), .ip2(n11630), .s(n11517), .op(
        n5727) );
  mux2_1 U13388 ( .ip1(\cache_data[8][81] ), .ip2(n11631), .s(n11517), .op(
        n5726) );
  mux2_1 U13389 ( .ip1(\cache_data[8][82] ), .ip2(n11632), .s(n11517), .op(
        n5725) );
  buf_1 U13390 ( .ip(n11517), .op(n11518) );
  mux2_1 U13391 ( .ip1(\cache_data[8][83] ), .ip2(n11633), .s(n11518), .op(
        n5724) );
  mux2_1 U13392 ( .ip1(\cache_data[8][84] ), .ip2(n11634), .s(n11518), .op(
        n5723) );
  mux2_1 U13393 ( .ip1(\cache_data[8][85] ), .ip2(n11635), .s(n11518), .op(
        n5722) );
  mux2_1 U13394 ( .ip1(\cache_data[8][86] ), .ip2(n11636), .s(n11518), .op(
        n5721) );
  mux2_1 U13395 ( .ip1(\cache_data[8][87] ), .ip2(n11637), .s(n11518), .op(
        n5720) );
  mux2_1 U13396 ( .ip1(\cache_data[8][88] ), .ip2(n11638), .s(n11517), .op(
        n5719) );
  mux2_1 U13397 ( .ip1(\cache_data[8][89] ), .ip2(n11640), .s(n11517), .op(
        n5718) );
  mux2_1 U13398 ( .ip1(\cache_data[8][90] ), .ip2(n11641), .s(n11518), .op(
        n5717) );
  mux2_1 U13399 ( .ip1(\cache_data[8][91] ), .ip2(n11642), .s(n11518), .op(
        n5716) );
  mux2_1 U13400 ( .ip1(\cache_data[8][92] ), .ip2(n11643), .s(n11518), .op(
        n5715) );
  mux2_1 U13401 ( .ip1(\cache_data[8][93] ), .ip2(n11644), .s(n11518), .op(
        n5714) );
  mux2_1 U13402 ( .ip1(\cache_data[8][94] ), .ip2(n11645), .s(n11518), .op(
        n5713) );
  mux2_1 U13403 ( .ip1(\cache_data[8][95] ), .ip2(n11647), .s(n11518), .op(
        n5712) );
  nor2_1 U13404 ( .ip1(n11613), .ip2(n8137), .op(n11519) );
  mux2_1 U13405 ( .ip1(\cache_data[8][96] ), .ip2(n11554), .s(n11519), .op(
        n5711) );
  mux2_1 U13406 ( .ip1(\cache_data[8][97] ), .ip2(n11555), .s(n11519), .op(
        n5710) );
  mux2_1 U13407 ( .ip1(\cache_data[8][98] ), .ip2(n11556), .s(n11519), .op(
        n5709) );
  mux2_1 U13408 ( .ip1(\cache_data[8][99] ), .ip2(n11557), .s(n11519), .op(
        n5708) );
  mux2_1 U13409 ( .ip1(\cache_data[8][100] ), .ip2(n11558), .s(n11519), .op(
        n5707) );
  mux2_1 U13410 ( .ip1(\cache_data[8][101] ), .ip2(n11559), .s(n11519), .op(
        n5706) );
  mux2_1 U13411 ( .ip1(\cache_data[8][102] ), .ip2(n11560), .s(n11519), .op(
        n5705) );
  mux2_1 U13412 ( .ip1(\cache_data[8][103] ), .ip2(n11561), .s(n11519), .op(
        n5704) );
  mux2_1 U13413 ( .ip1(\cache_data[8][104] ), .ip2(n11562), .s(n11519), .op(
        n5703) );
  mux2_1 U13414 ( .ip1(\cache_data[8][105] ), .ip2(n11563), .s(n11519), .op(
        n5702) );
  mux2_1 U13415 ( .ip1(\cache_data[8][106] ), .ip2(n11564), .s(n11519), .op(
        n5701) );
  mux2_1 U13416 ( .ip1(\cache_data[8][107] ), .ip2(n11565), .s(n11519), .op(
        n5700) );
  mux2_1 U13417 ( .ip1(\cache_data[8][108] ), .ip2(n11566), .s(n11519), .op(
        n5699) );
  mux2_1 U13418 ( .ip1(\cache_data[8][109] ), .ip2(n11567), .s(n11519), .op(
        n5698) );
  mux2_1 U13419 ( .ip1(\cache_data[8][110] ), .ip2(n11568), .s(n11519), .op(
        n5697) );
  mux2_1 U13420 ( .ip1(\cache_data[8][111] ), .ip2(n11569), .s(n11519), .op(
        n5696) );
  mux2_1 U13421 ( .ip1(\cache_data[8][112] ), .ip2(n11570), .s(n11519), .op(
        n5695) );
  mux2_1 U13422 ( .ip1(\cache_data[8][113] ), .ip2(n11571), .s(n11519), .op(
        n5694) );
  mux2_1 U13423 ( .ip1(\cache_data[8][114] ), .ip2(n11572), .s(n11519), .op(
        n5693) );
  buf_1 U13424 ( .ip(n11519), .op(n11520) );
  mux2_1 U13425 ( .ip1(\cache_data[8][115] ), .ip2(n11573), .s(n11520), .op(
        n5692) );
  mux2_1 U13426 ( .ip1(\cache_data[8][116] ), .ip2(n11574), .s(n11520), .op(
        n5691) );
  mux2_1 U13427 ( .ip1(\cache_data[8][117] ), .ip2(n11575), .s(n11520), .op(
        n5690) );
  mux2_1 U13428 ( .ip1(\cache_data[8][118] ), .ip2(n11576), .s(n11520), .op(
        n5689) );
  mux2_1 U13429 ( .ip1(\cache_data[8][119] ), .ip2(n11577), .s(n11520), .op(
        n5688) );
  mux2_1 U13430 ( .ip1(\cache_data[8][120] ), .ip2(n11578), .s(n11519), .op(
        n5687) );
  mux2_1 U13431 ( .ip1(\cache_data[8][121] ), .ip2(n11580), .s(n11519), .op(
        n5686) );
  mux2_1 U13432 ( .ip1(\cache_data[8][122] ), .ip2(n11581), .s(n11520), .op(
        n5685) );
  mux2_1 U13433 ( .ip1(\cache_data[8][123] ), .ip2(n11582), .s(n11520), .op(
        n5684) );
  mux2_1 U13434 ( .ip1(\cache_data[8][124] ), .ip2(n11583), .s(n11520), .op(
        n5683) );
  mux2_1 U13435 ( .ip1(\cache_data[8][125] ), .ip2(n11584), .s(n11520), .op(
        n5682) );
  mux2_1 U13436 ( .ip1(\cache_data[8][126] ), .ip2(n11585), .s(n11520), .op(
        n5681) );
  mux2_1 U13437 ( .ip1(\cache_data[8][127] ), .ip2(n11587), .s(n11520), .op(
        n5680) );
  nor2_1 U13438 ( .ip1(n11603), .ip2(n8144), .op(n11521) );
  mux2_1 U13439 ( .ip1(\cache_data[9][0] ), .ip2(n11614), .s(n11521), .op(
        n5679) );
  mux2_1 U13440 ( .ip1(\cache_data[9][1] ), .ip2(n11615), .s(n11521), .op(
        n5678) );
  mux2_1 U13441 ( .ip1(\cache_data[9][2] ), .ip2(n11616), .s(n11521), .op(
        n5677) );
  mux2_1 U13442 ( .ip1(\cache_data[9][3] ), .ip2(n11617), .s(n11521), .op(
        n5676) );
  mux2_1 U13443 ( .ip1(\cache_data[9][4] ), .ip2(n11618), .s(n11521), .op(
        n5675) );
  mux2_1 U13444 ( .ip1(\cache_data[9][5] ), .ip2(n11619), .s(n11521), .op(
        n5674) );
  mux2_1 U13445 ( .ip1(\cache_data[9][6] ), .ip2(n11620), .s(n11521), .op(
        n5673) );
  mux2_1 U13446 ( .ip1(\cache_data[9][7] ), .ip2(n11621), .s(n11521), .op(
        n5672) );
  mux2_1 U13447 ( .ip1(\cache_data[9][8] ), .ip2(n11622), .s(n11521), .op(
        n5671) );
  mux2_1 U13448 ( .ip1(\cache_data[9][9] ), .ip2(n11623), .s(n11521), .op(
        n5670) );
  mux2_1 U13449 ( .ip1(\cache_data[9][10] ), .ip2(n11624), .s(n11521), .op(
        n5669) );
  mux2_1 U13450 ( .ip1(\cache_data[9][11] ), .ip2(n11625), .s(n11521), .op(
        n5668) );
  mux2_1 U13451 ( .ip1(\cache_data[9][12] ), .ip2(n11626), .s(n11521), .op(
        n5667) );
  mux2_1 U13452 ( .ip1(\cache_data[9][13] ), .ip2(n11627), .s(n11521), .op(
        n5666) );
  mux2_1 U13453 ( .ip1(\cache_data[9][14] ), .ip2(n11628), .s(n11521), .op(
        n5665) );
  mux2_1 U13454 ( .ip1(\cache_data[9][15] ), .ip2(n11629), .s(n11521), .op(
        n5664) );
  mux2_1 U13455 ( .ip1(\cache_data[9][16] ), .ip2(n11630), .s(n11521), .op(
        n5663) );
  mux2_1 U13456 ( .ip1(\cache_data[9][17] ), .ip2(n11631), .s(n11521), .op(
        n5662) );
  mux2_1 U13457 ( .ip1(\cache_data[9][18] ), .ip2(n11632), .s(n11521), .op(
        n5661) );
  buf_1 U13458 ( .ip(n11521), .op(n11522) );
  mux2_1 U13459 ( .ip1(\cache_data[9][19] ), .ip2(n11633), .s(n11522), .op(
        n5660) );
  mux2_1 U13460 ( .ip1(\cache_data[9][20] ), .ip2(n11634), .s(n11522), .op(
        n5659) );
  mux2_1 U13461 ( .ip1(\cache_data[9][21] ), .ip2(n11635), .s(n11522), .op(
        n5658) );
  mux2_1 U13462 ( .ip1(\cache_data[9][22] ), .ip2(n11636), .s(n11522), .op(
        n5657) );
  mux2_1 U13463 ( .ip1(\cache_data[9][23] ), .ip2(n11637), .s(n11522), .op(
        n5656) );
  mux2_1 U13464 ( .ip1(\cache_data[9][24] ), .ip2(n11638), .s(n11521), .op(
        n5655) );
  mux2_1 U13465 ( .ip1(\cache_data[9][25] ), .ip2(n11640), .s(n11521), .op(
        n5654) );
  mux2_1 U13466 ( .ip1(\cache_data[9][26] ), .ip2(n11641), .s(n11522), .op(
        n5653) );
  mux2_1 U13467 ( .ip1(\cache_data[9][27] ), .ip2(n11642), .s(n11522), .op(
        n5652) );
  mux2_1 U13468 ( .ip1(\cache_data[9][28] ), .ip2(n11643), .s(n11522), .op(
        n5651) );
  mux2_1 U13469 ( .ip1(\cache_data[9][29] ), .ip2(n11644), .s(n11522), .op(
        n5650) );
  mux2_1 U13470 ( .ip1(\cache_data[9][30] ), .ip2(n11645), .s(n11522), .op(
        n5649) );
  mux2_1 U13471 ( .ip1(\cache_data[9][31] ), .ip2(n11647), .s(n11522), .op(
        n5648) );
  nor2_1 U13472 ( .ip1(n11606), .ip2(n8144), .op(n11523) );
  mux2_1 U13473 ( .ip1(\cache_data[9][32] ), .ip2(n11554), .s(n11523), .op(
        n5647) );
  mux2_1 U13474 ( .ip1(\cache_data[9][33] ), .ip2(n11555), .s(n11523), .op(
        n5646) );
  mux2_1 U13475 ( .ip1(\cache_data[9][34] ), .ip2(n11556), .s(n11523), .op(
        n5645) );
  mux2_1 U13476 ( .ip1(\cache_data[9][35] ), .ip2(n11557), .s(n11523), .op(
        n5644) );
  mux2_1 U13477 ( .ip1(\cache_data[9][36] ), .ip2(n11558), .s(n11523), .op(
        n5643) );
  mux2_1 U13478 ( .ip1(\cache_data[9][37] ), .ip2(n11559), .s(n11523), .op(
        n5642) );
  mux2_1 U13479 ( .ip1(\cache_data[9][38] ), .ip2(n11560), .s(n11523), .op(
        n5641) );
  mux2_1 U13480 ( .ip1(\cache_data[9][39] ), .ip2(n11561), .s(n11523), .op(
        n5640) );
  mux2_1 U13481 ( .ip1(\cache_data[9][40] ), .ip2(n11562), .s(n11523), .op(
        n5639) );
  mux2_1 U13482 ( .ip1(\cache_data[9][41] ), .ip2(n11563), .s(n11523), .op(
        n5638) );
  mux2_1 U13483 ( .ip1(\cache_data[9][42] ), .ip2(n11564), .s(n11523), .op(
        n5637) );
  mux2_1 U13484 ( .ip1(\cache_data[9][43] ), .ip2(n11565), .s(n11523), .op(
        n5636) );
  mux2_1 U13485 ( .ip1(\cache_data[9][44] ), .ip2(n11566), .s(n11523), .op(
        n5635) );
  mux2_1 U13486 ( .ip1(\cache_data[9][45] ), .ip2(n11567), .s(n11523), .op(
        n5634) );
  mux2_1 U13487 ( .ip1(\cache_data[9][46] ), .ip2(n11568), .s(n11523), .op(
        n5633) );
  mux2_1 U13488 ( .ip1(\cache_data[9][47] ), .ip2(n11569), .s(n11523), .op(
        n5632) );
  mux2_1 U13489 ( .ip1(\cache_data[9][48] ), .ip2(n11570), .s(n11523), .op(
        n5631) );
  mux2_1 U13490 ( .ip1(\cache_data[9][49] ), .ip2(n11571), .s(n11523), .op(
        n5630) );
  mux2_1 U13491 ( .ip1(\cache_data[9][50] ), .ip2(n11572), .s(n11523), .op(
        n5629) );
  buf_1 U13492 ( .ip(n11523), .op(n11524) );
  mux2_1 U13493 ( .ip1(\cache_data[9][51] ), .ip2(n11573), .s(n11524), .op(
        n5628) );
  mux2_1 U13494 ( .ip1(\cache_data[9][52] ), .ip2(n11574), .s(n11524), .op(
        n5627) );
  mux2_1 U13495 ( .ip1(\cache_data[9][53] ), .ip2(n11575), .s(n11524), .op(
        n5626) );
  mux2_1 U13496 ( .ip1(\cache_data[9][54] ), .ip2(n11576), .s(n11524), .op(
        n5625) );
  mux2_1 U13497 ( .ip1(\cache_data[9][55] ), .ip2(n11577), .s(n11524), .op(
        n5624) );
  mux2_1 U13498 ( .ip1(\cache_data[9][56] ), .ip2(n11578), .s(n11523), .op(
        n5623) );
  mux2_1 U13499 ( .ip1(\cache_data[9][57] ), .ip2(n11580), .s(n11523), .op(
        n5622) );
  mux2_1 U13500 ( .ip1(\cache_data[9][58] ), .ip2(n11581), .s(n11524), .op(
        n5621) );
  mux2_1 U13501 ( .ip1(\cache_data[9][59] ), .ip2(n11582), .s(n11524), .op(
        n5620) );
  mux2_1 U13502 ( .ip1(\cache_data[9][60] ), .ip2(n11583), .s(n11524), .op(
        n5619) );
  mux2_1 U13503 ( .ip1(\cache_data[9][61] ), .ip2(n11584), .s(n11524), .op(
        n5618) );
  mux2_1 U13504 ( .ip1(\cache_data[9][62] ), .ip2(n11585), .s(n11524), .op(
        n5617) );
  mux2_1 U13505 ( .ip1(\cache_data[9][63] ), .ip2(n11587), .s(n11524), .op(
        n5616) );
  nor2_1 U13506 ( .ip1(n11609), .ip2(n8144), .op(n11525) );
  mux2_1 U13507 ( .ip1(\cache_data[9][64] ), .ip2(n11614), .s(n11525), .op(
        n5615) );
  mux2_1 U13508 ( .ip1(\cache_data[9][65] ), .ip2(n11615), .s(n11525), .op(
        n5614) );
  mux2_1 U13509 ( .ip1(\cache_data[9][66] ), .ip2(n11616), .s(n11525), .op(
        n5613) );
  mux2_1 U13510 ( .ip1(\cache_data[9][67] ), .ip2(n11617), .s(n11525), .op(
        n5612) );
  mux2_1 U13511 ( .ip1(\cache_data[9][68] ), .ip2(n11618), .s(n11525), .op(
        n5611) );
  mux2_1 U13512 ( .ip1(\cache_data[9][69] ), .ip2(n11619), .s(n11525), .op(
        n5610) );
  mux2_1 U13513 ( .ip1(\cache_data[9][70] ), .ip2(n11620), .s(n11525), .op(
        n5609) );
  mux2_1 U13514 ( .ip1(\cache_data[9][71] ), .ip2(n11621), .s(n11525), .op(
        n5608) );
  mux2_1 U13515 ( .ip1(\cache_data[9][72] ), .ip2(n11622), .s(n11525), .op(
        n5607) );
  mux2_1 U13516 ( .ip1(\cache_data[9][73] ), .ip2(n11623), .s(n11525), .op(
        n5606) );
  mux2_1 U13517 ( .ip1(\cache_data[9][74] ), .ip2(n11624), .s(n11525), .op(
        n5605) );
  mux2_1 U13518 ( .ip1(\cache_data[9][75] ), .ip2(n11625), .s(n11525), .op(
        n5604) );
  mux2_1 U13519 ( .ip1(\cache_data[9][76] ), .ip2(n11626), .s(n11525), .op(
        n5603) );
  mux2_1 U13520 ( .ip1(\cache_data[9][77] ), .ip2(n11627), .s(n11525), .op(
        n5602) );
  mux2_1 U13521 ( .ip1(\cache_data[9][78] ), .ip2(n11628), .s(n11525), .op(
        n5601) );
  mux2_1 U13522 ( .ip1(\cache_data[9][79] ), .ip2(n11629), .s(n11525), .op(
        n5600) );
  mux2_1 U13523 ( .ip1(\cache_data[9][80] ), .ip2(n11630), .s(n11525), .op(
        n5599) );
  mux2_1 U13524 ( .ip1(\cache_data[9][81] ), .ip2(n11631), .s(n11525), .op(
        n5598) );
  mux2_1 U13525 ( .ip1(\cache_data[9][82] ), .ip2(n11632), .s(n11525), .op(
        n5597) );
  buf_1 U13526 ( .ip(n11525), .op(n11526) );
  mux2_1 U13527 ( .ip1(\cache_data[9][83] ), .ip2(n11633), .s(n11526), .op(
        n5596) );
  mux2_1 U13528 ( .ip1(\cache_data[9][84] ), .ip2(n11634), .s(n11526), .op(
        n5595) );
  mux2_1 U13529 ( .ip1(\cache_data[9][85] ), .ip2(n11635), .s(n11526), .op(
        n5594) );
  mux2_1 U13530 ( .ip1(\cache_data[9][86] ), .ip2(n11636), .s(n11526), .op(
        n5593) );
  mux2_1 U13531 ( .ip1(\cache_data[9][87] ), .ip2(n11637), .s(n11526), .op(
        n5592) );
  mux2_1 U13532 ( .ip1(\cache_data[9][88] ), .ip2(n11638), .s(n11525), .op(
        n5591) );
  mux2_1 U13533 ( .ip1(\cache_data[9][89] ), .ip2(n11640), .s(n11525), .op(
        n5590) );
  mux2_1 U13534 ( .ip1(\cache_data[9][90] ), .ip2(n11641), .s(n11526), .op(
        n5589) );
  mux2_1 U13535 ( .ip1(\cache_data[9][91] ), .ip2(n11642), .s(n11526), .op(
        n5588) );
  mux2_1 U13536 ( .ip1(\cache_data[9][92] ), .ip2(n11643), .s(n11526), .op(
        n5587) );
  mux2_1 U13537 ( .ip1(\cache_data[9][93] ), .ip2(n11644), .s(n11526), .op(
        n5586) );
  mux2_1 U13538 ( .ip1(\cache_data[9][94] ), .ip2(n11645), .s(n11526), .op(
        n5585) );
  mux2_1 U13539 ( .ip1(\cache_data[9][95] ), .ip2(n11647), .s(n11526), .op(
        n5584) );
  nor2_1 U13540 ( .ip1(n11613), .ip2(n8144), .op(n11527) );
  mux2_1 U13541 ( .ip1(\cache_data[9][96] ), .ip2(n11614), .s(n11527), .op(
        n5583) );
  mux2_1 U13542 ( .ip1(\cache_data[9][97] ), .ip2(n11615), .s(n11527), .op(
        n5582) );
  mux2_1 U13543 ( .ip1(\cache_data[9][98] ), .ip2(n11616), .s(n11527), .op(
        n5581) );
  mux2_1 U13544 ( .ip1(\cache_data[9][99] ), .ip2(n11617), .s(n11527), .op(
        n5580) );
  mux2_1 U13545 ( .ip1(\cache_data[9][100] ), .ip2(n11618), .s(n11527), .op(
        n5579) );
  mux2_1 U13546 ( .ip1(\cache_data[9][101] ), .ip2(n11619), .s(n11527), .op(
        n5578) );
  mux2_1 U13547 ( .ip1(\cache_data[9][102] ), .ip2(n11620), .s(n11527), .op(
        n5577) );
  mux2_1 U13548 ( .ip1(\cache_data[9][103] ), .ip2(n11621), .s(n11527), .op(
        n5576) );
  mux2_1 U13549 ( .ip1(\cache_data[9][104] ), .ip2(n11622), .s(n11527), .op(
        n5575) );
  mux2_1 U13550 ( .ip1(\cache_data[9][105] ), .ip2(n11623), .s(n11527), .op(
        n5574) );
  mux2_1 U13551 ( .ip1(\cache_data[9][106] ), .ip2(n11624), .s(n11527), .op(
        n5573) );
  mux2_1 U13552 ( .ip1(\cache_data[9][107] ), .ip2(n11625), .s(n11527), .op(
        n5572) );
  mux2_1 U13553 ( .ip1(\cache_data[9][108] ), .ip2(n11626), .s(n11527), .op(
        n5571) );
  mux2_1 U13554 ( .ip1(\cache_data[9][109] ), .ip2(n11627), .s(n11527), .op(
        n5570) );
  mux2_1 U13555 ( .ip1(\cache_data[9][110] ), .ip2(n11628), .s(n11527), .op(
        n5569) );
  mux2_1 U13556 ( .ip1(\cache_data[9][111] ), .ip2(n11629), .s(n11527), .op(
        n5568) );
  mux2_1 U13557 ( .ip1(\cache_data[9][112] ), .ip2(n11630), .s(n11527), .op(
        n5567) );
  mux2_1 U13558 ( .ip1(\cache_data[9][113] ), .ip2(n11631), .s(n11527), .op(
        n5566) );
  mux2_1 U13559 ( .ip1(\cache_data[9][114] ), .ip2(n11632), .s(n11527), .op(
        n5565) );
  buf_1 U13560 ( .ip(n11527), .op(n11528) );
  mux2_1 U13561 ( .ip1(\cache_data[9][115] ), .ip2(n11633), .s(n11528), .op(
        n5564) );
  mux2_1 U13562 ( .ip1(\cache_data[9][116] ), .ip2(n11634), .s(n11528), .op(
        n5563) );
  mux2_1 U13563 ( .ip1(\cache_data[9][117] ), .ip2(n11635), .s(n11528), .op(
        n5562) );
  mux2_1 U13564 ( .ip1(\cache_data[9][118] ), .ip2(n11636), .s(n11528), .op(
        n5561) );
  mux2_1 U13565 ( .ip1(\cache_data[9][119] ), .ip2(n11637), .s(n11528), .op(
        n5560) );
  mux2_1 U13566 ( .ip1(\cache_data[9][120] ), .ip2(n11638), .s(n11527), .op(
        n5559) );
  mux2_1 U13567 ( .ip1(\cache_data[9][121] ), .ip2(n11640), .s(n11527), .op(
        n5558) );
  mux2_1 U13568 ( .ip1(\cache_data[9][122] ), .ip2(n11641), .s(n11528), .op(
        n5557) );
  mux2_1 U13569 ( .ip1(\cache_data[9][123] ), .ip2(n11642), .s(n11528), .op(
        n5556) );
  mux2_1 U13570 ( .ip1(\cache_data[9][124] ), .ip2(n11643), .s(n11528), .op(
        n5555) );
  mux2_1 U13571 ( .ip1(\cache_data[9][125] ), .ip2(n11644), .s(n11528), .op(
        n5554) );
  mux2_1 U13572 ( .ip1(\cache_data[9][126] ), .ip2(n11645), .s(n11528), .op(
        n5553) );
  mux2_1 U13573 ( .ip1(\cache_data[9][127] ), .ip2(n11647), .s(n11528), .op(
        n5552) );
  nor2_1 U13574 ( .ip1(n11603), .ip2(n8146), .op(n11529) );
  mux2_1 U13575 ( .ip1(\cache_data[10][0] ), .ip2(n11554), .s(n11529), .op(
        n5551) );
  mux2_1 U13576 ( .ip1(\cache_data[10][1] ), .ip2(n11555), .s(n11529), .op(
        n5550) );
  mux2_1 U13577 ( .ip1(\cache_data[10][2] ), .ip2(n11556), .s(n11529), .op(
        n5549) );
  mux2_1 U13578 ( .ip1(\cache_data[10][3] ), .ip2(n11557), .s(n11529), .op(
        n5548) );
  mux2_1 U13579 ( .ip1(\cache_data[10][4] ), .ip2(n11558), .s(n11529), .op(
        n5547) );
  mux2_1 U13580 ( .ip1(\cache_data[10][5] ), .ip2(n11559), .s(n11529), .op(
        n5546) );
  mux2_1 U13581 ( .ip1(\cache_data[10][6] ), .ip2(n11560), .s(n11529), .op(
        n5545) );
  mux2_1 U13582 ( .ip1(\cache_data[10][7] ), .ip2(n11561), .s(n11529), .op(
        n5544) );
  mux2_1 U13583 ( .ip1(\cache_data[10][8] ), .ip2(n11562), .s(n11529), .op(
        n5543) );
  mux2_1 U13584 ( .ip1(\cache_data[10][9] ), .ip2(n11563), .s(n11529), .op(
        n5542) );
  mux2_1 U13585 ( .ip1(\cache_data[10][10] ), .ip2(n11564), .s(n11529), .op(
        n5541) );
  mux2_1 U13586 ( .ip1(\cache_data[10][11] ), .ip2(n11565), .s(n11529), .op(
        n5540) );
  mux2_1 U13587 ( .ip1(\cache_data[10][12] ), .ip2(n11566), .s(n11529), .op(
        n5539) );
  mux2_1 U13588 ( .ip1(\cache_data[10][13] ), .ip2(n11567), .s(n11529), .op(
        n5538) );
  mux2_1 U13589 ( .ip1(\cache_data[10][14] ), .ip2(n11568), .s(n11529), .op(
        n5537) );
  mux2_1 U13590 ( .ip1(\cache_data[10][15] ), .ip2(n11569), .s(n11529), .op(
        n5536) );
  mux2_1 U13591 ( .ip1(\cache_data[10][16] ), .ip2(n11570), .s(n11529), .op(
        n5535) );
  mux2_1 U13592 ( .ip1(\cache_data[10][17] ), .ip2(n11571), .s(n11529), .op(
        n5534) );
  mux2_1 U13593 ( .ip1(\cache_data[10][18] ), .ip2(n11572), .s(n11529), .op(
        n5533) );
  buf_1 U13594 ( .ip(n11529), .op(n11530) );
  mux2_1 U13595 ( .ip1(\cache_data[10][19] ), .ip2(n11573), .s(n11530), .op(
        n5532) );
  mux2_1 U13596 ( .ip1(\cache_data[10][20] ), .ip2(n11574), .s(n11530), .op(
        n5531) );
  mux2_1 U13597 ( .ip1(\cache_data[10][21] ), .ip2(n11575), .s(n11530), .op(
        n5530) );
  mux2_1 U13598 ( .ip1(\cache_data[10][22] ), .ip2(n11576), .s(n11530), .op(
        n5529) );
  mux2_1 U13599 ( .ip1(\cache_data[10][23] ), .ip2(n11577), .s(n11530), .op(
        n5528) );
  mux2_1 U13600 ( .ip1(\cache_data[10][24] ), .ip2(n11578), .s(n11529), .op(
        n5527) );
  mux2_1 U13601 ( .ip1(\cache_data[10][25] ), .ip2(n11580), .s(n11529), .op(
        n5526) );
  mux2_1 U13602 ( .ip1(\cache_data[10][26] ), .ip2(n11581), .s(n11530), .op(
        n5525) );
  mux2_1 U13603 ( .ip1(\cache_data[10][27] ), .ip2(n11582), .s(n11530), .op(
        n5524) );
  mux2_1 U13604 ( .ip1(\cache_data[10][28] ), .ip2(n11583), .s(n11530), .op(
        n5523) );
  mux2_1 U13605 ( .ip1(\cache_data[10][29] ), .ip2(n11584), .s(n11530), .op(
        n5522) );
  mux2_1 U13606 ( .ip1(\cache_data[10][30] ), .ip2(n11585), .s(n11530), .op(
        n5521) );
  mux2_1 U13607 ( .ip1(\cache_data[10][31] ), .ip2(n11587), .s(n11530), .op(
        n5520) );
  nor2_1 U13608 ( .ip1(n11606), .ip2(n8146), .op(n11531) );
  mux2_1 U13609 ( .ip1(\cache_data[10][32] ), .ip2(n11554), .s(n11531), .op(
        n5519) );
  mux2_1 U13610 ( .ip1(\cache_data[10][33] ), .ip2(n11555), .s(n11531), .op(
        n5518) );
  mux2_1 U13611 ( .ip1(\cache_data[10][34] ), .ip2(n11556), .s(n11531), .op(
        n5517) );
  mux2_1 U13612 ( .ip1(\cache_data[10][35] ), .ip2(n11557), .s(n11531), .op(
        n5516) );
  mux2_1 U13613 ( .ip1(\cache_data[10][36] ), .ip2(n11558), .s(n11531), .op(
        n5515) );
  mux2_1 U13614 ( .ip1(\cache_data[10][37] ), .ip2(n11559), .s(n11531), .op(
        n5514) );
  mux2_1 U13615 ( .ip1(\cache_data[10][38] ), .ip2(n11560), .s(n11531), .op(
        n5513) );
  mux2_1 U13616 ( .ip1(\cache_data[10][39] ), .ip2(n11561), .s(n11531), .op(
        n5512) );
  mux2_1 U13617 ( .ip1(\cache_data[10][40] ), .ip2(n11562), .s(n11531), .op(
        n5511) );
  mux2_1 U13618 ( .ip1(\cache_data[10][41] ), .ip2(n11563), .s(n11531), .op(
        n5510) );
  mux2_1 U13619 ( .ip1(\cache_data[10][42] ), .ip2(n11564), .s(n11531), .op(
        n5509) );
  mux2_1 U13620 ( .ip1(\cache_data[10][43] ), .ip2(n11565), .s(n11531), .op(
        n5508) );
  mux2_1 U13621 ( .ip1(\cache_data[10][44] ), .ip2(n11566), .s(n11531), .op(
        n5507) );
  mux2_1 U13622 ( .ip1(\cache_data[10][45] ), .ip2(n11567), .s(n11531), .op(
        n5506) );
  mux2_1 U13623 ( .ip1(\cache_data[10][46] ), .ip2(n11568), .s(n11531), .op(
        n5505) );
  mux2_1 U13624 ( .ip1(\cache_data[10][47] ), .ip2(n11569), .s(n11531), .op(
        n5504) );
  mux2_1 U13625 ( .ip1(\cache_data[10][48] ), .ip2(n11570), .s(n11531), .op(
        n5503) );
  mux2_1 U13626 ( .ip1(\cache_data[10][49] ), .ip2(n11571), .s(n11531), .op(
        n5502) );
  mux2_1 U13627 ( .ip1(\cache_data[10][50] ), .ip2(n11572), .s(n11531), .op(
        n5501) );
  buf_1 U13628 ( .ip(n11531), .op(n11532) );
  mux2_1 U13629 ( .ip1(\cache_data[10][51] ), .ip2(n11573), .s(n11532), .op(
        n5500) );
  mux2_1 U13630 ( .ip1(\cache_data[10][52] ), .ip2(n11574), .s(n11532), .op(
        n5499) );
  mux2_1 U13631 ( .ip1(\cache_data[10][53] ), .ip2(n11575), .s(n11532), .op(
        n5498) );
  mux2_1 U13632 ( .ip1(\cache_data[10][54] ), .ip2(n11576), .s(n11532), .op(
        n5497) );
  mux2_1 U13633 ( .ip1(\cache_data[10][55] ), .ip2(n11577), .s(n11532), .op(
        n5496) );
  mux2_1 U13634 ( .ip1(\cache_data[10][56] ), .ip2(n11578), .s(n11531), .op(
        n5495) );
  mux2_1 U13635 ( .ip1(\cache_data[10][57] ), .ip2(n11580), .s(n11531), .op(
        n5494) );
  mux2_1 U13636 ( .ip1(\cache_data[10][58] ), .ip2(n11581), .s(n11532), .op(
        n5493) );
  mux2_1 U13637 ( .ip1(\cache_data[10][59] ), .ip2(n11582), .s(n11532), .op(
        n5492) );
  mux2_1 U13638 ( .ip1(\cache_data[10][60] ), .ip2(n11583), .s(n11532), .op(
        n5491) );
  mux2_1 U13639 ( .ip1(\cache_data[10][61] ), .ip2(n11584), .s(n11532), .op(
        n5490) );
  mux2_1 U13640 ( .ip1(\cache_data[10][62] ), .ip2(n11585), .s(n11532), .op(
        n5489) );
  mux2_1 U13641 ( .ip1(\cache_data[10][63] ), .ip2(n11587), .s(n11532), .op(
        n5488) );
  nor2_1 U13642 ( .ip1(n11609), .ip2(n8146), .op(n11533) );
  mux2_1 U13643 ( .ip1(\cache_data[10][64] ), .ip2(n11554), .s(n11533), .op(
        n5487) );
  mux2_1 U13644 ( .ip1(\cache_data[10][65] ), .ip2(n11555), .s(n11533), .op(
        n5486) );
  mux2_1 U13645 ( .ip1(\cache_data[10][66] ), .ip2(n11556), .s(n11533), .op(
        n5485) );
  mux2_1 U13646 ( .ip1(\cache_data[10][67] ), .ip2(n11557), .s(n11533), .op(
        n5484) );
  mux2_1 U13647 ( .ip1(\cache_data[10][68] ), .ip2(n11558), .s(n11533), .op(
        n5483) );
  mux2_1 U13648 ( .ip1(\cache_data[10][69] ), .ip2(n11559), .s(n11533), .op(
        n5482) );
  mux2_1 U13649 ( .ip1(\cache_data[10][70] ), .ip2(n11560), .s(n11533), .op(
        n5481) );
  mux2_1 U13650 ( .ip1(\cache_data[10][71] ), .ip2(n11561), .s(n11533), .op(
        n5480) );
  mux2_1 U13651 ( .ip1(\cache_data[10][72] ), .ip2(n11562), .s(n11533), .op(
        n5479) );
  mux2_1 U13652 ( .ip1(\cache_data[10][73] ), .ip2(n11563), .s(n11533), .op(
        n5478) );
  mux2_1 U13653 ( .ip1(\cache_data[10][74] ), .ip2(n11564), .s(n11533), .op(
        n5477) );
  mux2_1 U13654 ( .ip1(\cache_data[10][75] ), .ip2(n11565), .s(n11533), .op(
        n5476) );
  mux2_1 U13655 ( .ip1(\cache_data[10][76] ), .ip2(n11566), .s(n11533), .op(
        n5475) );
  mux2_1 U13656 ( .ip1(\cache_data[10][77] ), .ip2(n11567), .s(n11533), .op(
        n5474) );
  mux2_1 U13657 ( .ip1(\cache_data[10][78] ), .ip2(n11568), .s(n11533), .op(
        n5473) );
  mux2_1 U13658 ( .ip1(\cache_data[10][79] ), .ip2(n11569), .s(n11533), .op(
        n5472) );
  mux2_1 U13659 ( .ip1(\cache_data[10][80] ), .ip2(n11570), .s(n11533), .op(
        n5471) );
  mux2_1 U13660 ( .ip1(\cache_data[10][81] ), .ip2(n11571), .s(n11533), .op(
        n5470) );
  mux2_1 U13661 ( .ip1(\cache_data[10][82] ), .ip2(n11572), .s(n11533), .op(
        n5469) );
  buf_1 U13662 ( .ip(n11533), .op(n11534) );
  mux2_1 U13663 ( .ip1(\cache_data[10][83] ), .ip2(n11573), .s(n11534), .op(
        n5468) );
  mux2_1 U13664 ( .ip1(\cache_data[10][84] ), .ip2(n11574), .s(n11534), .op(
        n5467) );
  mux2_1 U13665 ( .ip1(\cache_data[10][85] ), .ip2(n11575), .s(n11534), .op(
        n5466) );
  mux2_1 U13666 ( .ip1(\cache_data[10][86] ), .ip2(n11576), .s(n11534), .op(
        n5465) );
  mux2_1 U13667 ( .ip1(\cache_data[10][87] ), .ip2(n11577), .s(n11534), .op(
        n5464) );
  mux2_1 U13668 ( .ip1(\cache_data[10][88] ), .ip2(n11578), .s(n11533), .op(
        n5463) );
  mux2_1 U13669 ( .ip1(\cache_data[10][89] ), .ip2(n11580), .s(n11533), .op(
        n5462) );
  mux2_1 U13670 ( .ip1(\cache_data[10][90] ), .ip2(n11581), .s(n11534), .op(
        n5461) );
  mux2_1 U13671 ( .ip1(\cache_data[10][91] ), .ip2(n11582), .s(n11534), .op(
        n5460) );
  mux2_1 U13672 ( .ip1(\cache_data[10][92] ), .ip2(n11583), .s(n11534), .op(
        n5459) );
  mux2_1 U13673 ( .ip1(\cache_data[10][93] ), .ip2(n11584), .s(n11534), .op(
        n5458) );
  mux2_1 U13674 ( .ip1(\cache_data[10][94] ), .ip2(n11585), .s(n11534), .op(
        n5457) );
  mux2_1 U13675 ( .ip1(\cache_data[10][95] ), .ip2(n11587), .s(n11534), .op(
        n5456) );
  nor2_1 U13676 ( .ip1(n11613), .ip2(n8146), .op(n11535) );
  mux2_1 U13677 ( .ip1(\cache_data[10][96] ), .ip2(n11614), .s(n11535), .op(
        n5455) );
  mux2_1 U13678 ( .ip1(\cache_data[10][97] ), .ip2(n11615), .s(n11535), .op(
        n5454) );
  mux2_1 U13679 ( .ip1(\cache_data[10][98] ), .ip2(n11616), .s(n11535), .op(
        n5453) );
  mux2_1 U13680 ( .ip1(\cache_data[10][99] ), .ip2(n11617), .s(n11535), .op(
        n5452) );
  mux2_1 U13681 ( .ip1(\cache_data[10][100] ), .ip2(n11618), .s(n11535), .op(
        n5451) );
  mux2_1 U13682 ( .ip1(\cache_data[10][101] ), .ip2(n11619), .s(n11535), .op(
        n5450) );
  mux2_1 U13683 ( .ip1(\cache_data[10][102] ), .ip2(n11620), .s(n11535), .op(
        n5449) );
  mux2_1 U13684 ( .ip1(\cache_data[10][103] ), .ip2(n11621), .s(n11535), .op(
        n5448) );
  mux2_1 U13685 ( .ip1(\cache_data[10][104] ), .ip2(n11622), .s(n11535), .op(
        n5447) );
  mux2_1 U13686 ( .ip1(\cache_data[10][105] ), .ip2(n11623), .s(n11535), .op(
        n5446) );
  mux2_1 U13687 ( .ip1(\cache_data[10][106] ), .ip2(n11624), .s(n11535), .op(
        n5445) );
  mux2_1 U13688 ( .ip1(\cache_data[10][107] ), .ip2(n11625), .s(n11535), .op(
        n5444) );
  mux2_1 U13689 ( .ip1(\cache_data[10][108] ), .ip2(n11626), .s(n11535), .op(
        n5443) );
  mux2_1 U13690 ( .ip1(\cache_data[10][109] ), .ip2(n11627), .s(n11535), .op(
        n5442) );
  mux2_1 U13691 ( .ip1(\cache_data[10][110] ), .ip2(n11628), .s(n11535), .op(
        n5441) );
  mux2_1 U13692 ( .ip1(\cache_data[10][111] ), .ip2(n11629), .s(n11535), .op(
        n5440) );
  mux2_1 U13693 ( .ip1(\cache_data[10][112] ), .ip2(n11630), .s(n11535), .op(
        n5439) );
  mux2_1 U13694 ( .ip1(\cache_data[10][113] ), .ip2(n11631), .s(n11535), .op(
        n5438) );
  mux2_1 U13695 ( .ip1(\cache_data[10][114] ), .ip2(n11632), .s(n11535), .op(
        n5437) );
  buf_1 U13696 ( .ip(n11535), .op(n11536) );
  mux2_1 U13697 ( .ip1(\cache_data[10][115] ), .ip2(n11633), .s(n11536), .op(
        n5436) );
  mux2_1 U13698 ( .ip1(\cache_data[10][116] ), .ip2(n11634), .s(n11536), .op(
        n5435) );
  mux2_1 U13699 ( .ip1(\cache_data[10][117] ), .ip2(n11635), .s(n11536), .op(
        n5434) );
  mux2_1 U13700 ( .ip1(\cache_data[10][118] ), .ip2(n11636), .s(n11536), .op(
        n5433) );
  mux2_1 U13701 ( .ip1(\cache_data[10][119] ), .ip2(n11637), .s(n11536), .op(
        n5432) );
  mux2_1 U13702 ( .ip1(\cache_data[10][120] ), .ip2(n11638), .s(n11535), .op(
        n5431) );
  mux2_1 U13703 ( .ip1(\cache_data[10][121] ), .ip2(n11640), .s(n11535), .op(
        n5430) );
  mux2_1 U13704 ( .ip1(\cache_data[10][122] ), .ip2(n11641), .s(n11536), .op(
        n5429) );
  mux2_1 U13705 ( .ip1(\cache_data[10][123] ), .ip2(n11642), .s(n11536), .op(
        n5428) );
  mux2_1 U13706 ( .ip1(\cache_data[10][124] ), .ip2(n11643), .s(n11536), .op(
        n5427) );
  mux2_1 U13707 ( .ip1(\cache_data[10][125] ), .ip2(n11644), .s(n11536), .op(
        n5426) );
  mux2_1 U13708 ( .ip1(\cache_data[10][126] ), .ip2(n11645), .s(n11536), .op(
        n5425) );
  mux2_1 U13709 ( .ip1(\cache_data[10][127] ), .ip2(n11647), .s(n11536), .op(
        n5424) );
  nor2_1 U13710 ( .ip1(n11603), .ip2(n8151), .op(n11537) );
  mux2_1 U13711 ( .ip1(\cache_data[11][0] ), .ip2(n11554), .s(n11537), .op(
        n5423) );
  mux2_1 U13712 ( .ip1(\cache_data[11][1] ), .ip2(n11555), .s(n11537), .op(
        n5422) );
  mux2_1 U13713 ( .ip1(\cache_data[11][2] ), .ip2(n11556), .s(n11537), .op(
        n5421) );
  mux2_1 U13714 ( .ip1(\cache_data[11][3] ), .ip2(n11557), .s(n11537), .op(
        n5420) );
  mux2_1 U13715 ( .ip1(\cache_data[11][4] ), .ip2(n11558), .s(n11537), .op(
        n5419) );
  mux2_1 U13716 ( .ip1(\cache_data[11][5] ), .ip2(n11559), .s(n11537), .op(
        n5418) );
  mux2_1 U13717 ( .ip1(\cache_data[11][6] ), .ip2(n11560), .s(n11537), .op(
        n5417) );
  mux2_1 U13718 ( .ip1(\cache_data[11][7] ), .ip2(n11561), .s(n11537), .op(
        n5416) );
  mux2_1 U13719 ( .ip1(\cache_data[11][8] ), .ip2(n11562), .s(n11537), .op(
        n5415) );
  mux2_1 U13720 ( .ip1(\cache_data[11][9] ), .ip2(n11563), .s(n11537), .op(
        n5414) );
  mux2_1 U13721 ( .ip1(\cache_data[11][10] ), .ip2(n11564), .s(n11537), .op(
        n5413) );
  mux2_1 U13722 ( .ip1(\cache_data[11][11] ), .ip2(n11565), .s(n11537), .op(
        n5412) );
  mux2_1 U13723 ( .ip1(\cache_data[11][12] ), .ip2(n11566), .s(n11537), .op(
        n5411) );
  mux2_1 U13724 ( .ip1(\cache_data[11][13] ), .ip2(n11567), .s(n11537), .op(
        n5410) );
  mux2_1 U13725 ( .ip1(\cache_data[11][14] ), .ip2(n11568), .s(n11537), .op(
        n5409) );
  mux2_1 U13726 ( .ip1(\cache_data[11][15] ), .ip2(n11569), .s(n11537), .op(
        n5408) );
  mux2_1 U13727 ( .ip1(\cache_data[11][16] ), .ip2(n11570), .s(n11537), .op(
        n5407) );
  mux2_1 U13728 ( .ip1(\cache_data[11][17] ), .ip2(n11571), .s(n11537), .op(
        n5406) );
  mux2_1 U13729 ( .ip1(\cache_data[11][18] ), .ip2(n11572), .s(n11537), .op(
        n5405) );
  buf_1 U13730 ( .ip(n11537), .op(n11538) );
  mux2_1 U13731 ( .ip1(\cache_data[11][19] ), .ip2(n11573), .s(n11538), .op(
        n5404) );
  mux2_1 U13732 ( .ip1(\cache_data[11][20] ), .ip2(n11574), .s(n11538), .op(
        n5403) );
  mux2_1 U13733 ( .ip1(\cache_data[11][21] ), .ip2(n11575), .s(n11538), .op(
        n5402) );
  mux2_1 U13734 ( .ip1(\cache_data[11][22] ), .ip2(n11576), .s(n11538), .op(
        n5401) );
  mux2_1 U13735 ( .ip1(\cache_data[11][23] ), .ip2(n11577), .s(n11538), .op(
        n5400) );
  mux2_1 U13736 ( .ip1(\cache_data[11][24] ), .ip2(n11578), .s(n11537), .op(
        n5399) );
  mux2_1 U13737 ( .ip1(\cache_data[11][25] ), .ip2(n11580), .s(n11537), .op(
        n5398) );
  mux2_1 U13738 ( .ip1(\cache_data[11][26] ), .ip2(n11581), .s(n11538), .op(
        n5397) );
  mux2_1 U13739 ( .ip1(\cache_data[11][27] ), .ip2(n11582), .s(n11538), .op(
        n5396) );
  mux2_1 U13740 ( .ip1(\cache_data[11][28] ), .ip2(n11583), .s(n11538), .op(
        n5395) );
  mux2_1 U13741 ( .ip1(\cache_data[11][29] ), .ip2(n11584), .s(n11538), .op(
        n5394) );
  mux2_1 U13742 ( .ip1(\cache_data[11][30] ), .ip2(n11585), .s(n11538), .op(
        n5393) );
  mux2_1 U13743 ( .ip1(\cache_data[11][31] ), .ip2(n11587), .s(n11538), .op(
        n5392) );
  nor2_1 U13744 ( .ip1(n11606), .ip2(n8151), .op(n11539) );
  mux2_1 U13745 ( .ip1(\cache_data[11][32] ), .ip2(n11554), .s(n11539), .op(
        n5391) );
  mux2_1 U13746 ( .ip1(\cache_data[11][33] ), .ip2(n11555), .s(n11539), .op(
        n5390) );
  mux2_1 U13747 ( .ip1(\cache_data[11][34] ), .ip2(n11556), .s(n11539), .op(
        n5389) );
  mux2_1 U13748 ( .ip1(\cache_data[11][35] ), .ip2(n11557), .s(n11539), .op(
        n5388) );
  mux2_1 U13749 ( .ip1(\cache_data[11][36] ), .ip2(n11558), .s(n11539), .op(
        n5387) );
  mux2_1 U13750 ( .ip1(\cache_data[11][37] ), .ip2(n11559), .s(n11539), .op(
        n5386) );
  mux2_1 U13751 ( .ip1(\cache_data[11][38] ), .ip2(n11560), .s(n11539), .op(
        n5385) );
  mux2_1 U13752 ( .ip1(\cache_data[11][39] ), .ip2(n11561), .s(n11539), .op(
        n5384) );
  mux2_1 U13753 ( .ip1(\cache_data[11][40] ), .ip2(n11562), .s(n11539), .op(
        n5383) );
  mux2_1 U13754 ( .ip1(\cache_data[11][41] ), .ip2(n11563), .s(n11539), .op(
        n5382) );
  mux2_1 U13755 ( .ip1(\cache_data[11][42] ), .ip2(n11564), .s(n11539), .op(
        n5381) );
  mux2_1 U13756 ( .ip1(\cache_data[11][43] ), .ip2(n11565), .s(n11539), .op(
        n5380) );
  mux2_1 U13757 ( .ip1(\cache_data[11][44] ), .ip2(n11566), .s(n11539), .op(
        n5379) );
  mux2_1 U13758 ( .ip1(\cache_data[11][45] ), .ip2(n11567), .s(n11539), .op(
        n5378) );
  mux2_1 U13759 ( .ip1(\cache_data[11][46] ), .ip2(n11568), .s(n11539), .op(
        n5377) );
  mux2_1 U13760 ( .ip1(\cache_data[11][47] ), .ip2(n11569), .s(n11539), .op(
        n5376) );
  mux2_1 U13761 ( .ip1(\cache_data[11][48] ), .ip2(n11570), .s(n11539), .op(
        n5375) );
  mux2_1 U13762 ( .ip1(\cache_data[11][49] ), .ip2(n11571), .s(n11539), .op(
        n5374) );
  mux2_1 U13763 ( .ip1(\cache_data[11][50] ), .ip2(n11572), .s(n11539), .op(
        n5373) );
  buf_1 U13764 ( .ip(n11539), .op(n11540) );
  mux2_1 U13765 ( .ip1(\cache_data[11][51] ), .ip2(n11573), .s(n11540), .op(
        n5372) );
  mux2_1 U13766 ( .ip1(\cache_data[11][52] ), .ip2(n11574), .s(n11540), .op(
        n5371) );
  mux2_1 U13767 ( .ip1(\cache_data[11][53] ), .ip2(n11575), .s(n11540), .op(
        n5370) );
  mux2_1 U13768 ( .ip1(\cache_data[11][54] ), .ip2(n11576), .s(n11540), .op(
        n5369) );
  mux2_1 U13769 ( .ip1(\cache_data[11][55] ), .ip2(n11577), .s(n11540), .op(
        n5368) );
  mux2_1 U13770 ( .ip1(\cache_data[11][56] ), .ip2(n11578), .s(n11539), .op(
        n5367) );
  mux2_1 U13771 ( .ip1(\cache_data[11][57] ), .ip2(n11580), .s(n11539), .op(
        n5366) );
  mux2_1 U13772 ( .ip1(\cache_data[11][58] ), .ip2(n11581), .s(n11540), .op(
        n5365) );
  mux2_1 U13773 ( .ip1(\cache_data[11][59] ), .ip2(n11582), .s(n11540), .op(
        n5364) );
  mux2_1 U13774 ( .ip1(\cache_data[11][60] ), .ip2(n11583), .s(n11540), .op(
        n5363) );
  mux2_1 U13775 ( .ip1(\cache_data[11][61] ), .ip2(n11584), .s(n11540), .op(
        n5362) );
  mux2_1 U13776 ( .ip1(\cache_data[11][62] ), .ip2(n11585), .s(n11540), .op(
        n5361) );
  mux2_1 U13777 ( .ip1(\cache_data[11][63] ), .ip2(n11587), .s(n11540), .op(
        n5360) );
  nor2_1 U13778 ( .ip1(n11609), .ip2(n8151), .op(n11541) );
  mux2_1 U13779 ( .ip1(\cache_data[11][64] ), .ip2(n11554), .s(n11541), .op(
        n5359) );
  mux2_1 U13780 ( .ip1(\cache_data[11][65] ), .ip2(n11555), .s(n11541), .op(
        n5358) );
  mux2_1 U13781 ( .ip1(\cache_data[11][66] ), .ip2(n11556), .s(n11541), .op(
        n5357) );
  mux2_1 U13782 ( .ip1(\cache_data[11][67] ), .ip2(n11557), .s(n11541), .op(
        n5356) );
  mux2_1 U13783 ( .ip1(\cache_data[11][68] ), .ip2(n11558), .s(n11541), .op(
        n5355) );
  mux2_1 U13784 ( .ip1(\cache_data[11][69] ), .ip2(n11559), .s(n11541), .op(
        n5354) );
  mux2_1 U13785 ( .ip1(\cache_data[11][70] ), .ip2(n11560), .s(n11541), .op(
        n5353) );
  mux2_1 U13786 ( .ip1(\cache_data[11][71] ), .ip2(n11561), .s(n11541), .op(
        n5352) );
  mux2_1 U13787 ( .ip1(\cache_data[11][72] ), .ip2(n11562), .s(n11541), .op(
        n5351) );
  mux2_1 U13788 ( .ip1(\cache_data[11][73] ), .ip2(n11563), .s(n11541), .op(
        n5350) );
  mux2_1 U13789 ( .ip1(\cache_data[11][74] ), .ip2(n11564), .s(n11541), .op(
        n5349) );
  mux2_1 U13790 ( .ip1(\cache_data[11][75] ), .ip2(n11565), .s(n11541), .op(
        n5348) );
  mux2_1 U13791 ( .ip1(\cache_data[11][76] ), .ip2(n11566), .s(n11541), .op(
        n5347) );
  mux2_1 U13792 ( .ip1(\cache_data[11][77] ), .ip2(n11567), .s(n11541), .op(
        n5346) );
  mux2_1 U13793 ( .ip1(\cache_data[11][78] ), .ip2(n11568), .s(n11541), .op(
        n5345) );
  mux2_1 U13794 ( .ip1(\cache_data[11][79] ), .ip2(n11569), .s(n11541), .op(
        n5344) );
  mux2_1 U13795 ( .ip1(\cache_data[11][80] ), .ip2(n11570), .s(n11541), .op(
        n5343) );
  mux2_1 U13796 ( .ip1(\cache_data[11][81] ), .ip2(n11571), .s(n11541), .op(
        n5342) );
  mux2_1 U13797 ( .ip1(\cache_data[11][82] ), .ip2(n11572), .s(n11541), .op(
        n5341) );
  buf_1 U13798 ( .ip(n11541), .op(n11542) );
  mux2_1 U13799 ( .ip1(\cache_data[11][83] ), .ip2(n11573), .s(n11542), .op(
        n5340) );
  mux2_1 U13800 ( .ip1(\cache_data[11][84] ), .ip2(n11574), .s(n11542), .op(
        n5339) );
  mux2_1 U13801 ( .ip1(\cache_data[11][85] ), .ip2(n11575), .s(n11542), .op(
        n5338) );
  mux2_1 U13802 ( .ip1(\cache_data[11][86] ), .ip2(n11576), .s(n11542), .op(
        n5337) );
  mux2_1 U13803 ( .ip1(\cache_data[11][87] ), .ip2(n11577), .s(n11542), .op(
        n5336) );
  mux2_1 U13804 ( .ip1(\cache_data[11][88] ), .ip2(n11578), .s(n11541), .op(
        n5335) );
  mux2_1 U13805 ( .ip1(\cache_data[11][89] ), .ip2(n11580), .s(n11541), .op(
        n5334) );
  mux2_1 U13806 ( .ip1(\cache_data[11][90] ), .ip2(n11581), .s(n11542), .op(
        n5333) );
  mux2_1 U13807 ( .ip1(\cache_data[11][91] ), .ip2(n11582), .s(n11542), .op(
        n5332) );
  mux2_1 U13808 ( .ip1(\cache_data[11][92] ), .ip2(n11583), .s(n11542), .op(
        n5331) );
  mux2_1 U13809 ( .ip1(\cache_data[11][93] ), .ip2(n11584), .s(n11542), .op(
        n5330) );
  mux2_1 U13810 ( .ip1(\cache_data[11][94] ), .ip2(n11585), .s(n11542), .op(
        n5329) );
  mux2_1 U13811 ( .ip1(\cache_data[11][95] ), .ip2(n11587), .s(n11542), .op(
        n5328) );
  nor2_1 U13812 ( .ip1(n11613), .ip2(n8151), .op(n11543) );
  mux2_1 U13813 ( .ip1(\cache_data[11][96] ), .ip2(n11614), .s(n11543), .op(
        n5327) );
  mux2_1 U13814 ( .ip1(\cache_data[11][97] ), .ip2(n11615), .s(n11543), .op(
        n5326) );
  mux2_1 U13815 ( .ip1(\cache_data[11][98] ), .ip2(n11616), .s(n11543), .op(
        n5325) );
  mux2_1 U13816 ( .ip1(\cache_data[11][99] ), .ip2(n11617), .s(n11543), .op(
        n5324) );
  mux2_1 U13817 ( .ip1(\cache_data[11][100] ), .ip2(n11618), .s(n11543), .op(
        n5323) );
  mux2_1 U13818 ( .ip1(\cache_data[11][101] ), .ip2(n11619), .s(n11543), .op(
        n5322) );
  mux2_1 U13819 ( .ip1(\cache_data[11][102] ), .ip2(n11620), .s(n11543), .op(
        n5321) );
  mux2_1 U13820 ( .ip1(\cache_data[11][103] ), .ip2(n11621), .s(n11543), .op(
        n5320) );
  mux2_1 U13821 ( .ip1(\cache_data[11][104] ), .ip2(n11622), .s(n11543), .op(
        n5319) );
  mux2_1 U13822 ( .ip1(\cache_data[11][105] ), .ip2(n11623), .s(n11543), .op(
        n5318) );
  mux2_1 U13823 ( .ip1(\cache_data[11][106] ), .ip2(n11624), .s(n11543), .op(
        n5317) );
  mux2_1 U13824 ( .ip1(\cache_data[11][107] ), .ip2(n11625), .s(n11543), .op(
        n5316) );
  mux2_1 U13825 ( .ip1(\cache_data[11][108] ), .ip2(n11626), .s(n11543), .op(
        n5315) );
  mux2_1 U13826 ( .ip1(\cache_data[11][109] ), .ip2(n11627), .s(n11543), .op(
        n5314) );
  mux2_1 U13827 ( .ip1(\cache_data[11][110] ), .ip2(n11628), .s(n11543), .op(
        n5313) );
  mux2_1 U13828 ( .ip1(\cache_data[11][111] ), .ip2(n11629), .s(n11543), .op(
        n5312) );
  mux2_1 U13829 ( .ip1(\cache_data[11][112] ), .ip2(n11630), .s(n11543), .op(
        n5311) );
  mux2_1 U13830 ( .ip1(\cache_data[11][113] ), .ip2(n11631), .s(n11543), .op(
        n5310) );
  mux2_1 U13831 ( .ip1(\cache_data[11][114] ), .ip2(n11632), .s(n11543), .op(
        n5309) );
  buf_1 U13832 ( .ip(n11543), .op(n11544) );
  mux2_1 U13833 ( .ip1(\cache_data[11][115] ), .ip2(n11633), .s(n11544), .op(
        n5308) );
  mux2_1 U13834 ( .ip1(\cache_data[11][116] ), .ip2(n11634), .s(n11544), .op(
        n5307) );
  mux2_1 U13835 ( .ip1(\cache_data[11][117] ), .ip2(n11635), .s(n11544), .op(
        n5306) );
  mux2_1 U13836 ( .ip1(\cache_data[11][118] ), .ip2(n11636), .s(n11544), .op(
        n5305) );
  mux2_1 U13837 ( .ip1(\cache_data[11][119] ), .ip2(n11637), .s(n11544), .op(
        n5304) );
  mux2_1 U13838 ( .ip1(\cache_data[11][120] ), .ip2(n11638), .s(n11543), .op(
        n5303) );
  mux2_1 U13839 ( .ip1(\cache_data[11][121] ), .ip2(n11640), .s(n11543), .op(
        n5302) );
  mux2_1 U13840 ( .ip1(\cache_data[11][122] ), .ip2(n11641), .s(n11544), .op(
        n5301) );
  mux2_1 U13841 ( .ip1(\cache_data[11][123] ), .ip2(n11642), .s(n11544), .op(
        n5300) );
  mux2_1 U13842 ( .ip1(\cache_data[11][124] ), .ip2(n11643), .s(n11544), .op(
        n5299) );
  mux2_1 U13843 ( .ip1(\cache_data[11][125] ), .ip2(n11644), .s(n11544), .op(
        n5298) );
  mux2_1 U13844 ( .ip1(\cache_data[11][126] ), .ip2(n11645), .s(n11544), .op(
        n5297) );
  mux2_1 U13845 ( .ip1(\cache_data[11][127] ), .ip2(n11647), .s(n11544), .op(
        n5296) );
  nor2_1 U13846 ( .ip1(n11603), .ip2(n11551), .op(n11545) );
  mux2_1 U13847 ( .ip1(\cache_data[12][0] ), .ip2(n11554), .s(n11545), .op(
        n5295) );
  mux2_1 U13848 ( .ip1(\cache_data[12][1] ), .ip2(n11555), .s(n11545), .op(
        n5294) );
  mux2_1 U13849 ( .ip1(\cache_data[12][2] ), .ip2(n11556), .s(n11545), .op(
        n5293) );
  mux2_1 U13850 ( .ip1(\cache_data[12][3] ), .ip2(n11557), .s(n11545), .op(
        n5292) );
  mux2_1 U13851 ( .ip1(\cache_data[12][4] ), .ip2(n11558), .s(n11545), .op(
        n5291) );
  mux2_1 U13852 ( .ip1(\cache_data[12][5] ), .ip2(n11559), .s(n11545), .op(
        n5290) );
  mux2_1 U13853 ( .ip1(\cache_data[12][6] ), .ip2(n11560), .s(n11545), .op(
        n5289) );
  mux2_1 U13854 ( .ip1(\cache_data[12][7] ), .ip2(n11561), .s(n11545), .op(
        n5288) );
  mux2_1 U13855 ( .ip1(\cache_data[12][8] ), .ip2(n11562), .s(n11545), .op(
        n5287) );
  mux2_1 U13856 ( .ip1(\cache_data[12][9] ), .ip2(n11563), .s(n11545), .op(
        n5286) );
  mux2_1 U13857 ( .ip1(\cache_data[12][10] ), .ip2(n11564), .s(n11545), .op(
        n5285) );
  mux2_1 U13858 ( .ip1(\cache_data[12][11] ), .ip2(n11565), .s(n11545), .op(
        n5284) );
  mux2_1 U13859 ( .ip1(\cache_data[12][12] ), .ip2(n11566), .s(n11545), .op(
        n5283) );
  mux2_1 U13860 ( .ip1(\cache_data[12][13] ), .ip2(n11567), .s(n11545), .op(
        n5282) );
  mux2_1 U13861 ( .ip1(\cache_data[12][14] ), .ip2(n11568), .s(n11545), .op(
        n5281) );
  mux2_1 U13862 ( .ip1(\cache_data[12][15] ), .ip2(n11569), .s(n11545), .op(
        n5280) );
  mux2_1 U13863 ( .ip1(\cache_data[12][16] ), .ip2(n11570), .s(n11545), .op(
        n5279) );
  mux2_1 U13864 ( .ip1(\cache_data[12][17] ), .ip2(n11571), .s(n11545), .op(
        n5278) );
  mux2_1 U13865 ( .ip1(\cache_data[12][18] ), .ip2(n11572), .s(n11545), .op(
        n5277) );
  buf_1 U13866 ( .ip(n11545), .op(n11546) );
  mux2_1 U13867 ( .ip1(\cache_data[12][19] ), .ip2(n11573), .s(n11546), .op(
        n5276) );
  mux2_1 U13868 ( .ip1(\cache_data[12][20] ), .ip2(n11574), .s(n11546), .op(
        n5275) );
  mux2_1 U13869 ( .ip1(\cache_data[12][21] ), .ip2(n11575), .s(n11546), .op(
        n5274) );
  mux2_1 U13870 ( .ip1(\cache_data[12][22] ), .ip2(n11576), .s(n11546), .op(
        n5273) );
  mux2_1 U13871 ( .ip1(\cache_data[12][23] ), .ip2(n11577), .s(n11546), .op(
        n5272) );
  mux2_1 U13872 ( .ip1(\cache_data[12][24] ), .ip2(n11578), .s(n11545), .op(
        n5271) );
  mux2_1 U13873 ( .ip1(\cache_data[12][25] ), .ip2(n11580), .s(n11545), .op(
        n5270) );
  mux2_1 U13874 ( .ip1(\cache_data[12][26] ), .ip2(n11581), .s(n11546), .op(
        n5269) );
  mux2_1 U13875 ( .ip1(\cache_data[12][27] ), .ip2(n11582), .s(n11546), .op(
        n5268) );
  mux2_1 U13876 ( .ip1(\cache_data[12][28] ), .ip2(n11583), .s(n11546), .op(
        n5267) );
  mux2_1 U13877 ( .ip1(\cache_data[12][29] ), .ip2(n11584), .s(n11546), .op(
        n5266) );
  mux2_1 U13878 ( .ip1(\cache_data[12][30] ), .ip2(n11585), .s(n11546), .op(
        n5265) );
  mux2_1 U13879 ( .ip1(\cache_data[12][31] ), .ip2(n11587), .s(n11546), .op(
        n5264) );
  nor2_1 U13880 ( .ip1(n11606), .ip2(n11551), .op(n11547) );
  mux2_1 U13881 ( .ip1(\cache_data[12][32] ), .ip2(n11554), .s(n11547), .op(
        n5263) );
  mux2_1 U13882 ( .ip1(\cache_data[12][33] ), .ip2(n11555), .s(n11547), .op(
        n5262) );
  mux2_1 U13883 ( .ip1(\cache_data[12][34] ), .ip2(n11556), .s(n11547), .op(
        n5261) );
  mux2_1 U13884 ( .ip1(\cache_data[12][35] ), .ip2(n11557), .s(n11547), .op(
        n5260) );
  mux2_1 U13885 ( .ip1(\cache_data[12][36] ), .ip2(n11558), .s(n11547), .op(
        n5259) );
  mux2_1 U13886 ( .ip1(\cache_data[12][37] ), .ip2(n11559), .s(n11547), .op(
        n5258) );
  mux2_1 U13887 ( .ip1(\cache_data[12][38] ), .ip2(n11560), .s(n11547), .op(
        n5257) );
  mux2_1 U13888 ( .ip1(\cache_data[12][39] ), .ip2(n11561), .s(n11547), .op(
        n5256) );
  mux2_1 U13889 ( .ip1(\cache_data[12][40] ), .ip2(n11562), .s(n11547), .op(
        n5255) );
  mux2_1 U13890 ( .ip1(\cache_data[12][41] ), .ip2(n11563), .s(n11547), .op(
        n5254) );
  mux2_1 U13891 ( .ip1(\cache_data[12][42] ), .ip2(n11564), .s(n11547), .op(
        n5253) );
  mux2_1 U13892 ( .ip1(\cache_data[12][43] ), .ip2(n11565), .s(n11547), .op(
        n5252) );
  mux2_1 U13893 ( .ip1(\cache_data[12][44] ), .ip2(n11566), .s(n11547), .op(
        n5251) );
  mux2_1 U13894 ( .ip1(\cache_data[12][45] ), .ip2(n11567), .s(n11547), .op(
        n5250) );
  mux2_1 U13895 ( .ip1(\cache_data[12][46] ), .ip2(n11568), .s(n11547), .op(
        n5249) );
  mux2_1 U13896 ( .ip1(\cache_data[12][47] ), .ip2(n11569), .s(n11547), .op(
        n5248) );
  mux2_1 U13897 ( .ip1(\cache_data[12][48] ), .ip2(n11570), .s(n11547), .op(
        n5247) );
  mux2_1 U13898 ( .ip1(\cache_data[12][49] ), .ip2(n11571), .s(n11547), .op(
        n5246) );
  mux2_1 U13899 ( .ip1(\cache_data[12][50] ), .ip2(n11572), .s(n11547), .op(
        n5245) );
  buf_1 U13900 ( .ip(n11547), .op(n11548) );
  mux2_1 U13901 ( .ip1(\cache_data[12][51] ), .ip2(n11573), .s(n11548), .op(
        n5244) );
  mux2_1 U13902 ( .ip1(\cache_data[12][52] ), .ip2(n11574), .s(n11548), .op(
        n5243) );
  mux2_1 U13903 ( .ip1(\cache_data[12][53] ), .ip2(n11575), .s(n11548), .op(
        n5242) );
  mux2_1 U13904 ( .ip1(\cache_data[12][54] ), .ip2(n11576), .s(n11548), .op(
        n5241) );
  mux2_1 U13905 ( .ip1(\cache_data[12][55] ), .ip2(n11577), .s(n11548), .op(
        n5240) );
  mux2_1 U13906 ( .ip1(\cache_data[12][56] ), .ip2(n11578), .s(n11547), .op(
        n5239) );
  mux2_1 U13907 ( .ip1(\cache_data[12][57] ), .ip2(n11580), .s(n11547), .op(
        n5238) );
  mux2_1 U13908 ( .ip1(\cache_data[12][58] ), .ip2(n11581), .s(n11548), .op(
        n5237) );
  mux2_1 U13909 ( .ip1(\cache_data[12][59] ), .ip2(n11582), .s(n11548), .op(
        n5236) );
  mux2_1 U13910 ( .ip1(\cache_data[12][60] ), .ip2(n11583), .s(n11548), .op(
        n5235) );
  mux2_1 U13911 ( .ip1(\cache_data[12][61] ), .ip2(n11584), .s(n11548), .op(
        n5234) );
  mux2_1 U13912 ( .ip1(\cache_data[12][62] ), .ip2(n11585), .s(n11548), .op(
        n5233) );
  mux2_1 U13913 ( .ip1(\cache_data[12][63] ), .ip2(n11587), .s(n11548), .op(
        n5232) );
  nor2_1 U13914 ( .ip1(n11609), .ip2(n11551), .op(n11549) );
  mux2_1 U13915 ( .ip1(\cache_data[12][64] ), .ip2(n11554), .s(n11549), .op(
        n5231) );
  mux2_1 U13916 ( .ip1(\cache_data[12][65] ), .ip2(n11555), .s(n11549), .op(
        n5230) );
  mux2_1 U13917 ( .ip1(\cache_data[12][66] ), .ip2(n11556), .s(n11549), .op(
        n5229) );
  mux2_1 U13918 ( .ip1(\cache_data[12][67] ), .ip2(n11557), .s(n11549), .op(
        n5228) );
  mux2_1 U13919 ( .ip1(\cache_data[12][68] ), .ip2(n11558), .s(n11549), .op(
        n5227) );
  mux2_1 U13920 ( .ip1(\cache_data[12][69] ), .ip2(n11559), .s(n11549), .op(
        n5226) );
  mux2_1 U13921 ( .ip1(\cache_data[12][70] ), .ip2(n11560), .s(n11549), .op(
        n5225) );
  mux2_1 U13922 ( .ip1(\cache_data[12][71] ), .ip2(n11561), .s(n11549), .op(
        n5224) );
  mux2_1 U13923 ( .ip1(\cache_data[12][72] ), .ip2(n11562), .s(n11549), .op(
        n5223) );
  mux2_1 U13924 ( .ip1(\cache_data[12][73] ), .ip2(n11563), .s(n11549), .op(
        n5222) );
  mux2_1 U13925 ( .ip1(\cache_data[12][74] ), .ip2(n11564), .s(n11549), .op(
        n5221) );
  mux2_1 U13926 ( .ip1(\cache_data[12][75] ), .ip2(n11565), .s(n11549), .op(
        n5220) );
  mux2_1 U13927 ( .ip1(\cache_data[12][76] ), .ip2(n11566), .s(n11549), .op(
        n5219) );
  mux2_1 U13928 ( .ip1(\cache_data[12][77] ), .ip2(n11567), .s(n11549), .op(
        n5218) );
  mux2_1 U13929 ( .ip1(\cache_data[12][78] ), .ip2(n11568), .s(n11549), .op(
        n5217) );
  mux2_1 U13930 ( .ip1(\cache_data[12][79] ), .ip2(n11569), .s(n11549), .op(
        n5216) );
  mux2_1 U13931 ( .ip1(\cache_data[12][80] ), .ip2(n11570), .s(n11549), .op(
        n5215) );
  mux2_1 U13932 ( .ip1(\cache_data[12][81] ), .ip2(n11571), .s(n11549), .op(
        n5214) );
  mux2_1 U13933 ( .ip1(\cache_data[12][82] ), .ip2(n11572), .s(n11549), .op(
        n5213) );
  buf_1 U13934 ( .ip(n11549), .op(n11550) );
  mux2_1 U13935 ( .ip1(\cache_data[12][83] ), .ip2(n11573), .s(n11550), .op(
        n5212) );
  mux2_1 U13936 ( .ip1(\cache_data[12][84] ), .ip2(n11574), .s(n11550), .op(
        n5211) );
  mux2_1 U13937 ( .ip1(\cache_data[12][85] ), .ip2(n11575), .s(n11550), .op(
        n5210) );
  mux2_1 U13938 ( .ip1(\cache_data[12][86] ), .ip2(n11576), .s(n11550), .op(
        n5209) );
  mux2_1 U13939 ( .ip1(\cache_data[12][87] ), .ip2(n11577), .s(n11550), .op(
        n5208) );
  mux2_1 U13940 ( .ip1(\cache_data[12][88] ), .ip2(n11578), .s(n11549), .op(
        n5207) );
  mux2_1 U13941 ( .ip1(\cache_data[12][89] ), .ip2(n11580), .s(n11549), .op(
        n5206) );
  mux2_1 U13942 ( .ip1(\cache_data[12][90] ), .ip2(n11581), .s(n11550), .op(
        n5205) );
  mux2_1 U13943 ( .ip1(\cache_data[12][91] ), .ip2(n11582), .s(n11550), .op(
        n5204) );
  mux2_1 U13944 ( .ip1(\cache_data[12][92] ), .ip2(n11583), .s(n11550), .op(
        n5203) );
  mux2_1 U13945 ( .ip1(\cache_data[12][93] ), .ip2(n11584), .s(n11550), .op(
        n5202) );
  mux2_1 U13946 ( .ip1(\cache_data[12][94] ), .ip2(n11585), .s(n11550), .op(
        n5201) );
  mux2_1 U13947 ( .ip1(\cache_data[12][95] ), .ip2(n11587), .s(n11550), .op(
        n5200) );
  nor2_1 U13948 ( .ip1(n11613), .ip2(n11551), .op(n11552) );
  mux2_1 U13949 ( .ip1(\cache_data[12][96] ), .ip2(n11554), .s(n11552), .op(
        n5199) );
  mux2_1 U13950 ( .ip1(\cache_data[12][97] ), .ip2(n11555), .s(n11552), .op(
        n5198) );
  mux2_1 U13951 ( .ip1(\cache_data[12][98] ), .ip2(n11556), .s(n11552), .op(
        n5197) );
  mux2_1 U13952 ( .ip1(\cache_data[12][99] ), .ip2(n11557), .s(n11552), .op(
        n5196) );
  mux2_1 U13953 ( .ip1(\cache_data[12][100] ), .ip2(n11558), .s(n11552), .op(
        n5195) );
  mux2_1 U13954 ( .ip1(\cache_data[12][101] ), .ip2(n11559), .s(n11552), .op(
        n5194) );
  mux2_1 U13955 ( .ip1(\cache_data[12][102] ), .ip2(n11560), .s(n11552), .op(
        n5193) );
  mux2_1 U13956 ( .ip1(\cache_data[12][103] ), .ip2(n11561), .s(n11552), .op(
        n5192) );
  mux2_1 U13957 ( .ip1(\cache_data[12][104] ), .ip2(n11562), .s(n11552), .op(
        n5191) );
  mux2_1 U13958 ( .ip1(\cache_data[12][105] ), .ip2(n11563), .s(n11552), .op(
        n5190) );
  mux2_1 U13959 ( .ip1(\cache_data[12][106] ), .ip2(n11564), .s(n11552), .op(
        n5189) );
  mux2_1 U13960 ( .ip1(\cache_data[12][107] ), .ip2(n11565), .s(n11552), .op(
        n5188) );
  mux2_1 U13961 ( .ip1(\cache_data[12][108] ), .ip2(n11566), .s(n11552), .op(
        n5187) );
  mux2_1 U13962 ( .ip1(\cache_data[12][109] ), .ip2(n11567), .s(n11552), .op(
        n5186) );
  mux2_1 U13963 ( .ip1(\cache_data[12][110] ), .ip2(n11568), .s(n11552), .op(
        n5185) );
  mux2_1 U13964 ( .ip1(\cache_data[12][111] ), .ip2(n11569), .s(n11552), .op(
        n5184) );
  mux2_1 U13965 ( .ip1(\cache_data[12][112] ), .ip2(n11570), .s(n11552), .op(
        n5183) );
  mux2_1 U13966 ( .ip1(\cache_data[12][113] ), .ip2(n11571), .s(n11552), .op(
        n5182) );
  mux2_1 U13967 ( .ip1(\cache_data[12][114] ), .ip2(n11572), .s(n11552), .op(
        n5181) );
  buf_1 U13968 ( .ip(n11552), .op(n11553) );
  mux2_1 U13969 ( .ip1(\cache_data[12][115] ), .ip2(n11573), .s(n11553), .op(
        n5180) );
  mux2_1 U13970 ( .ip1(\cache_data[12][116] ), .ip2(n11574), .s(n11553), .op(
        n5179) );
  mux2_1 U13971 ( .ip1(\cache_data[12][117] ), .ip2(n11575), .s(n11553), .op(
        n5178) );
  mux2_1 U13972 ( .ip1(\cache_data[12][118] ), .ip2(n11576), .s(n11553), .op(
        n5177) );
  mux2_1 U13973 ( .ip1(\cache_data[12][119] ), .ip2(n11577), .s(n11553), .op(
        n5176) );
  mux2_1 U13974 ( .ip1(\cache_data[12][120] ), .ip2(n11578), .s(n11552), .op(
        n5175) );
  mux2_1 U13975 ( .ip1(\cache_data[12][121] ), .ip2(n11580), .s(n11552), .op(
        n5174) );
  mux2_1 U13976 ( .ip1(\cache_data[12][122] ), .ip2(n11581), .s(n11553), .op(
        n5173) );
  mux2_1 U13977 ( .ip1(\cache_data[12][123] ), .ip2(n11582), .s(n11553), .op(
        n5172) );
  mux2_1 U13978 ( .ip1(\cache_data[12][124] ), .ip2(n11583), .s(n11553), .op(
        n5171) );
  mux2_1 U13979 ( .ip1(\cache_data[12][125] ), .ip2(n11584), .s(n11553), .op(
        n5170) );
  mux2_1 U13980 ( .ip1(\cache_data[12][126] ), .ip2(n11585), .s(n11553), .op(
        n5169) );
  mux2_1 U13981 ( .ip1(\cache_data[12][127] ), .ip2(n11587), .s(n11553), .op(
        n5168) );
  nor2_1 U13982 ( .ip1(n11603), .ip2(n8145), .op(n11579) );
  mux2_1 U13983 ( .ip1(\cache_data[13][0] ), .ip2(n11554), .s(n11579), .op(
        n5167) );
  mux2_1 U13984 ( .ip1(\cache_data[13][1] ), .ip2(n11555), .s(n11579), .op(
        n5166) );
  mux2_1 U13985 ( .ip1(\cache_data[13][2] ), .ip2(n11556), .s(n11579), .op(
        n5165) );
  mux2_1 U13986 ( .ip1(\cache_data[13][3] ), .ip2(n11557), .s(n11579), .op(
        n5164) );
  mux2_1 U13987 ( .ip1(\cache_data[13][4] ), .ip2(n11558), .s(n11579), .op(
        n5163) );
  mux2_1 U13988 ( .ip1(\cache_data[13][5] ), .ip2(n11559), .s(n11579), .op(
        n5162) );
  mux2_1 U13989 ( .ip1(\cache_data[13][6] ), .ip2(n11560), .s(n11579), .op(
        n5161) );
  mux2_1 U13990 ( .ip1(\cache_data[13][7] ), .ip2(n11561), .s(n11579), .op(
        n5160) );
  mux2_1 U13991 ( .ip1(\cache_data[13][8] ), .ip2(n11562), .s(n11579), .op(
        n5159) );
  mux2_1 U13992 ( .ip1(\cache_data[13][9] ), .ip2(n11563), .s(n11579), .op(
        n5158) );
  mux2_1 U13993 ( .ip1(\cache_data[13][10] ), .ip2(n11564), .s(n11579), .op(
        n5157) );
  mux2_1 U13994 ( .ip1(\cache_data[13][11] ), .ip2(n11565), .s(n11579), .op(
        n5156) );
  mux2_1 U13995 ( .ip1(\cache_data[13][12] ), .ip2(n11566), .s(n11579), .op(
        n5155) );
  mux2_1 U13996 ( .ip1(\cache_data[13][13] ), .ip2(n11567), .s(n11579), .op(
        n5154) );
  mux2_1 U13997 ( .ip1(\cache_data[13][14] ), .ip2(n11568), .s(n11579), .op(
        n5153) );
  mux2_1 U13998 ( .ip1(\cache_data[13][15] ), .ip2(n11569), .s(n11579), .op(
        n5152) );
  mux2_1 U13999 ( .ip1(\cache_data[13][16] ), .ip2(n11570), .s(n11579), .op(
        n5151) );
  mux2_1 U14000 ( .ip1(\cache_data[13][17] ), .ip2(n11571), .s(n11579), .op(
        n5150) );
  mux2_1 U14001 ( .ip1(\cache_data[13][18] ), .ip2(n11572), .s(n11579), .op(
        n5149) );
  buf_1 U14002 ( .ip(n11579), .op(n11586) );
  mux2_1 U14003 ( .ip1(\cache_data[13][19] ), .ip2(n11573), .s(n11586), .op(
        n5148) );
  mux2_1 U14004 ( .ip1(\cache_data[13][20] ), .ip2(n11574), .s(n11586), .op(
        n5147) );
  mux2_1 U14005 ( .ip1(\cache_data[13][21] ), .ip2(n11575), .s(n11586), .op(
        n5146) );
  mux2_1 U14006 ( .ip1(\cache_data[13][22] ), .ip2(n11576), .s(n11586), .op(
        n5145) );
  mux2_1 U14007 ( .ip1(\cache_data[13][23] ), .ip2(n11577), .s(n11586), .op(
        n5144) );
  mux2_1 U14008 ( .ip1(\cache_data[13][24] ), .ip2(n11578), .s(n11579), .op(
        n5143) );
  mux2_1 U14009 ( .ip1(\cache_data[13][25] ), .ip2(n11580), .s(n11579), .op(
        n5142) );
  mux2_1 U14010 ( .ip1(\cache_data[13][26] ), .ip2(n11581), .s(n11586), .op(
        n5141) );
  mux2_1 U14011 ( .ip1(\cache_data[13][27] ), .ip2(n11582), .s(n11586), .op(
        n5140) );
  mux2_1 U14012 ( .ip1(\cache_data[13][28] ), .ip2(n11583), .s(n11586), .op(
        n5139) );
  mux2_1 U14013 ( .ip1(\cache_data[13][29] ), .ip2(n11584), .s(n11586), .op(
        n5138) );
  mux2_1 U14014 ( .ip1(\cache_data[13][30] ), .ip2(n11585), .s(n11586), .op(
        n5137) );
  mux2_1 U14015 ( .ip1(\cache_data[13][31] ), .ip2(n11587), .s(n11586), .op(
        n5136) );
  nor2_1 U14016 ( .ip1(n11606), .ip2(n8145), .op(n11588) );
  mux2_1 U14017 ( .ip1(\cache_data[13][32] ), .ip2(n11614), .s(n11588), .op(
        n5135) );
  mux2_1 U14018 ( .ip1(\cache_data[13][33] ), .ip2(n11615), .s(n11588), .op(
        n5134) );
  mux2_1 U14019 ( .ip1(\cache_data[13][34] ), .ip2(n11616), .s(n11588), .op(
        n5133) );
  mux2_1 U14020 ( .ip1(\cache_data[13][35] ), .ip2(n11617), .s(n11588), .op(
        n5132) );
  mux2_1 U14021 ( .ip1(\cache_data[13][36] ), .ip2(n11618), .s(n11588), .op(
        n5131) );
  mux2_1 U14022 ( .ip1(\cache_data[13][37] ), .ip2(n11619), .s(n11588), .op(
        n5130) );
  mux2_1 U14023 ( .ip1(\cache_data[13][38] ), .ip2(n11620), .s(n11588), .op(
        n5129) );
  mux2_1 U14024 ( .ip1(\cache_data[13][39] ), .ip2(n11621), .s(n11588), .op(
        n5128) );
  mux2_1 U14025 ( .ip1(\cache_data[13][40] ), .ip2(n11622), .s(n11588), .op(
        n5127) );
  mux2_1 U14026 ( .ip1(\cache_data[13][41] ), .ip2(n11623), .s(n11588), .op(
        n5126) );
  mux2_1 U14027 ( .ip1(\cache_data[13][42] ), .ip2(n11624), .s(n11588), .op(
        n5125) );
  mux2_1 U14028 ( .ip1(\cache_data[13][43] ), .ip2(n11625), .s(n11588), .op(
        n5124) );
  mux2_1 U14029 ( .ip1(\cache_data[13][44] ), .ip2(n11626), .s(n11588), .op(
        n5123) );
  mux2_1 U14030 ( .ip1(\cache_data[13][45] ), .ip2(n11627), .s(n11588), .op(
        n5122) );
  mux2_1 U14031 ( .ip1(\cache_data[13][46] ), .ip2(n11628), .s(n11588), .op(
        n5121) );
  mux2_1 U14032 ( .ip1(\cache_data[13][47] ), .ip2(n11629), .s(n11588), .op(
        n5120) );
  mux2_1 U14033 ( .ip1(\cache_data[13][48] ), .ip2(n11630), .s(n11588), .op(
        n5119) );
  mux2_1 U14034 ( .ip1(\cache_data[13][49] ), .ip2(n11631), .s(n11588), .op(
        n5118) );
  mux2_1 U14035 ( .ip1(\cache_data[13][50] ), .ip2(n11632), .s(n11588), .op(
        n5117) );
  buf_1 U14036 ( .ip(n11588), .op(n11589) );
  mux2_1 U14037 ( .ip1(\cache_data[13][51] ), .ip2(n11633), .s(n11589), .op(
        n5116) );
  mux2_1 U14038 ( .ip1(\cache_data[13][52] ), .ip2(n11634), .s(n11589), .op(
        n5115) );
  mux2_1 U14039 ( .ip1(\cache_data[13][53] ), .ip2(n11635), .s(n11589), .op(
        n5114) );
  mux2_1 U14040 ( .ip1(\cache_data[13][54] ), .ip2(n11636), .s(n11589), .op(
        n5113) );
  mux2_1 U14041 ( .ip1(\cache_data[13][55] ), .ip2(n11637), .s(n11589), .op(
        n5112) );
  mux2_1 U14042 ( .ip1(\cache_data[13][56] ), .ip2(n11638), .s(n11588), .op(
        n5111) );
  mux2_1 U14043 ( .ip1(\cache_data[13][57] ), .ip2(n11640), .s(n11588), .op(
        n5110) );
  mux2_1 U14044 ( .ip1(\cache_data[13][58] ), .ip2(n11641), .s(n11589), .op(
        n5109) );
  mux2_1 U14045 ( .ip1(\cache_data[13][59] ), .ip2(n11642), .s(n11589), .op(
        n5108) );
  mux2_1 U14046 ( .ip1(\cache_data[13][60] ), .ip2(n11643), .s(n11589), .op(
        n5107) );
  mux2_1 U14047 ( .ip1(\cache_data[13][61] ), .ip2(n11644), .s(n11589), .op(
        n5106) );
  mux2_1 U14048 ( .ip1(\cache_data[13][62] ), .ip2(n11645), .s(n11589), .op(
        n5105) );
  mux2_1 U14049 ( .ip1(\cache_data[13][63] ), .ip2(n11647), .s(n11589), .op(
        n5104) );
  nor2_1 U14050 ( .ip1(n11609), .ip2(n8145), .op(n11590) );
  mux2_1 U14051 ( .ip1(\cache_data[13][64] ), .ip2(n11614), .s(n11590), .op(
        n5103) );
  mux2_1 U14052 ( .ip1(\cache_data[13][65] ), .ip2(n11615), .s(n11590), .op(
        n5102) );
  mux2_1 U14053 ( .ip1(\cache_data[13][66] ), .ip2(n11616), .s(n11590), .op(
        n5101) );
  mux2_1 U14054 ( .ip1(\cache_data[13][67] ), .ip2(n11617), .s(n11590), .op(
        n5100) );
  mux2_1 U14055 ( .ip1(\cache_data[13][68] ), .ip2(n11618), .s(n11590), .op(
        n5099) );
  mux2_1 U14056 ( .ip1(\cache_data[13][69] ), .ip2(n11619), .s(n11590), .op(
        n5098) );
  mux2_1 U14057 ( .ip1(\cache_data[13][70] ), .ip2(n11620), .s(n11590), .op(
        n5097) );
  mux2_1 U14058 ( .ip1(\cache_data[13][71] ), .ip2(n11621), .s(n11590), .op(
        n5096) );
  mux2_1 U14059 ( .ip1(\cache_data[13][72] ), .ip2(n11622), .s(n11590), .op(
        n5095) );
  mux2_1 U14060 ( .ip1(\cache_data[13][73] ), .ip2(n11623), .s(n11590), .op(
        n5094) );
  mux2_1 U14061 ( .ip1(\cache_data[13][74] ), .ip2(n11624), .s(n11590), .op(
        n5093) );
  mux2_1 U14062 ( .ip1(\cache_data[13][75] ), .ip2(n11625), .s(n11590), .op(
        n5092) );
  mux2_1 U14063 ( .ip1(\cache_data[13][76] ), .ip2(n11626), .s(n11590), .op(
        n5091) );
  mux2_1 U14064 ( .ip1(\cache_data[13][77] ), .ip2(n11627), .s(n11590), .op(
        n5090) );
  mux2_1 U14065 ( .ip1(\cache_data[13][78] ), .ip2(n11628), .s(n11590), .op(
        n5089) );
  mux2_1 U14066 ( .ip1(\cache_data[13][79] ), .ip2(n11629), .s(n11590), .op(
        n5088) );
  mux2_1 U14067 ( .ip1(\cache_data[13][80] ), .ip2(n11630), .s(n11590), .op(
        n5087) );
  mux2_1 U14068 ( .ip1(\cache_data[13][81] ), .ip2(n11631), .s(n11590), .op(
        n5086) );
  mux2_1 U14069 ( .ip1(\cache_data[13][82] ), .ip2(n11632), .s(n11590), .op(
        n5085) );
  buf_1 U14070 ( .ip(n11590), .op(n11591) );
  mux2_1 U14071 ( .ip1(\cache_data[13][83] ), .ip2(n11633), .s(n11591), .op(
        n5084) );
  mux2_1 U14072 ( .ip1(\cache_data[13][84] ), .ip2(n11634), .s(n11591), .op(
        n5083) );
  mux2_1 U14073 ( .ip1(\cache_data[13][85] ), .ip2(n11635), .s(n11591), .op(
        n5082) );
  mux2_1 U14074 ( .ip1(\cache_data[13][86] ), .ip2(n11636), .s(n11591), .op(
        n5081) );
  mux2_1 U14075 ( .ip1(\cache_data[13][87] ), .ip2(n11637), .s(n11591), .op(
        n5080) );
  mux2_1 U14076 ( .ip1(\cache_data[13][88] ), .ip2(n11638), .s(n11590), .op(
        n5079) );
  mux2_1 U14077 ( .ip1(\cache_data[13][89] ), .ip2(n11640), .s(n11590), .op(
        n5078) );
  mux2_1 U14078 ( .ip1(\cache_data[13][90] ), .ip2(n11641), .s(n11591), .op(
        n5077) );
  mux2_1 U14079 ( .ip1(\cache_data[13][91] ), .ip2(n11642), .s(n11591), .op(
        n5076) );
  mux2_1 U14080 ( .ip1(\cache_data[13][92] ), .ip2(n11643), .s(n11591), .op(
        n5075) );
  mux2_1 U14081 ( .ip1(\cache_data[13][93] ), .ip2(n11644), .s(n11591), .op(
        n5074) );
  mux2_1 U14082 ( .ip1(\cache_data[13][94] ), .ip2(n11645), .s(n11591), .op(
        n5073) );
  mux2_1 U14083 ( .ip1(\cache_data[13][95] ), .ip2(n11647), .s(n11591), .op(
        n5072) );
  nor2_1 U14084 ( .ip1(n11613), .ip2(n8145), .op(n11592) );
  mux2_1 U14085 ( .ip1(\cache_data[13][96] ), .ip2(n11614), .s(n11592), .op(
        n5071) );
  mux2_1 U14086 ( .ip1(\cache_data[13][97] ), .ip2(n11615), .s(n11592), .op(
        n5070) );
  mux2_1 U14087 ( .ip1(\cache_data[13][98] ), .ip2(n11616), .s(n11592), .op(
        n5069) );
  mux2_1 U14088 ( .ip1(\cache_data[13][99] ), .ip2(n11617), .s(n11592), .op(
        n5068) );
  mux2_1 U14089 ( .ip1(\cache_data[13][100] ), .ip2(n11618), .s(n11592), .op(
        n5067) );
  mux2_1 U14090 ( .ip1(\cache_data[13][101] ), .ip2(n11619), .s(n11592), .op(
        n5066) );
  mux2_1 U14091 ( .ip1(\cache_data[13][102] ), .ip2(n11620), .s(n11592), .op(
        n5065) );
  mux2_1 U14092 ( .ip1(\cache_data[13][103] ), .ip2(n11621), .s(n11592), .op(
        n5064) );
  mux2_1 U14093 ( .ip1(\cache_data[13][104] ), .ip2(n11622), .s(n11592), .op(
        n5063) );
  mux2_1 U14094 ( .ip1(\cache_data[13][105] ), .ip2(n11623), .s(n11592), .op(
        n5062) );
  mux2_1 U14095 ( .ip1(\cache_data[13][106] ), .ip2(n11624), .s(n11592), .op(
        n5061) );
  mux2_1 U14096 ( .ip1(\cache_data[13][107] ), .ip2(n11625), .s(n11592), .op(
        n5060) );
  mux2_1 U14097 ( .ip1(\cache_data[13][108] ), .ip2(n11626), .s(n11592), .op(
        n5059) );
  mux2_1 U14098 ( .ip1(\cache_data[13][109] ), .ip2(n11627), .s(n11592), .op(
        n5058) );
  mux2_1 U14099 ( .ip1(\cache_data[13][110] ), .ip2(n11628), .s(n11592), .op(
        n5057) );
  mux2_1 U14100 ( .ip1(\cache_data[13][111] ), .ip2(n11629), .s(n11592), .op(
        n5056) );
  mux2_1 U14101 ( .ip1(\cache_data[13][112] ), .ip2(n11630), .s(n11592), .op(
        n5055) );
  mux2_1 U14102 ( .ip1(\cache_data[13][113] ), .ip2(n11631), .s(n11592), .op(
        n5054) );
  mux2_1 U14103 ( .ip1(\cache_data[13][114] ), .ip2(n11632), .s(n11592), .op(
        n5053) );
  buf_1 U14104 ( .ip(n11592), .op(n11593) );
  mux2_1 U14105 ( .ip1(\cache_data[13][115] ), .ip2(n11633), .s(n11593), .op(
        n5052) );
  mux2_1 U14106 ( .ip1(\cache_data[13][116] ), .ip2(n11634), .s(n11593), .op(
        n5051) );
  mux2_1 U14107 ( .ip1(\cache_data[13][117] ), .ip2(n11635), .s(n11593), .op(
        n5050) );
  mux2_1 U14108 ( .ip1(\cache_data[13][118] ), .ip2(n11636), .s(n11593), .op(
        n5049) );
  mux2_1 U14109 ( .ip1(\cache_data[13][119] ), .ip2(n11637), .s(n11593), .op(
        n5048) );
  mux2_1 U14110 ( .ip1(\cache_data[13][120] ), .ip2(n11638), .s(n11592), .op(
        n5047) );
  mux2_1 U14111 ( .ip1(\cache_data[13][121] ), .ip2(n11640), .s(n11592), .op(
        n5046) );
  mux2_1 U14112 ( .ip1(\cache_data[13][122] ), .ip2(n11641), .s(n11593), .op(
        n5045) );
  mux2_1 U14113 ( .ip1(\cache_data[13][123] ), .ip2(n11642), .s(n11593), .op(
        n5044) );
  mux2_1 U14114 ( .ip1(\cache_data[13][124] ), .ip2(n11643), .s(n11593), .op(
        n5043) );
  mux2_1 U14115 ( .ip1(\cache_data[13][125] ), .ip2(n11644), .s(n11593), .op(
        n5042) );
  mux2_1 U14116 ( .ip1(\cache_data[13][126] ), .ip2(n11645), .s(n11593), .op(
        n5041) );
  mux2_1 U14117 ( .ip1(\cache_data[13][127] ), .ip2(n11647), .s(n11593), .op(
        n5040) );
  nor2_1 U14118 ( .ip1(n11603), .ip2(n11600), .op(n11594) );
  mux2_1 U14119 ( .ip1(\cache_data[14][0] ), .ip2(n11614), .s(n11594), .op(
        n5039) );
  mux2_1 U14120 ( .ip1(\cache_data[14][1] ), .ip2(n11615), .s(n11594), .op(
        n5038) );
  mux2_1 U14121 ( .ip1(\cache_data[14][2] ), .ip2(n11616), .s(n11594), .op(
        n5037) );
  mux2_1 U14122 ( .ip1(\cache_data[14][3] ), .ip2(n11617), .s(n11594), .op(
        n5036) );
  mux2_1 U14123 ( .ip1(\cache_data[14][4] ), .ip2(n11618), .s(n11594), .op(
        n5035) );
  mux2_1 U14124 ( .ip1(\cache_data[14][5] ), .ip2(n11619), .s(n11594), .op(
        n5034) );
  mux2_1 U14125 ( .ip1(\cache_data[14][6] ), .ip2(n11620), .s(n11594), .op(
        n5033) );
  mux2_1 U14126 ( .ip1(\cache_data[14][7] ), .ip2(n11621), .s(n11594), .op(
        n5032) );
  mux2_1 U14127 ( .ip1(\cache_data[14][8] ), .ip2(n11622), .s(n11594), .op(
        n5031) );
  mux2_1 U14128 ( .ip1(\cache_data[14][9] ), .ip2(n11623), .s(n11594), .op(
        n5030) );
  mux2_1 U14129 ( .ip1(\cache_data[14][10] ), .ip2(n11624), .s(n11594), .op(
        n5029) );
  mux2_1 U14130 ( .ip1(\cache_data[14][11] ), .ip2(n11625), .s(n11594), .op(
        n5028) );
  mux2_1 U14131 ( .ip1(\cache_data[14][12] ), .ip2(n11626), .s(n11594), .op(
        n5027) );
  mux2_1 U14132 ( .ip1(\cache_data[14][13] ), .ip2(n11627), .s(n11594), .op(
        n5026) );
  mux2_1 U14133 ( .ip1(\cache_data[14][14] ), .ip2(n11628), .s(n11594), .op(
        n5025) );
  mux2_1 U14134 ( .ip1(\cache_data[14][15] ), .ip2(n11629), .s(n11594), .op(
        n5024) );
  mux2_1 U14135 ( .ip1(\cache_data[14][16] ), .ip2(n11630), .s(n11594), .op(
        n5023) );
  mux2_1 U14136 ( .ip1(\cache_data[14][17] ), .ip2(n11631), .s(n11594), .op(
        n5022) );
  mux2_1 U14137 ( .ip1(\cache_data[14][18] ), .ip2(n11632), .s(n11594), .op(
        n5021) );
  buf_1 U14138 ( .ip(n11594), .op(n11595) );
  mux2_1 U14139 ( .ip1(\cache_data[14][19] ), .ip2(n11633), .s(n11595), .op(
        n5020) );
  mux2_1 U14140 ( .ip1(\cache_data[14][20] ), .ip2(n11634), .s(n11595), .op(
        n5019) );
  mux2_1 U14141 ( .ip1(\cache_data[14][21] ), .ip2(n11635), .s(n11595), .op(
        n5018) );
  mux2_1 U14142 ( .ip1(\cache_data[14][22] ), .ip2(n11636), .s(n11595), .op(
        n5017) );
  mux2_1 U14143 ( .ip1(\cache_data[14][23] ), .ip2(n11637), .s(n11595), .op(
        n5016) );
  mux2_1 U14144 ( .ip1(\cache_data[14][24] ), .ip2(n11638), .s(n11594), .op(
        n5015) );
  mux2_1 U14145 ( .ip1(\cache_data[14][25] ), .ip2(n11640), .s(n11594), .op(
        n5014) );
  mux2_1 U14146 ( .ip1(\cache_data[14][26] ), .ip2(n11641), .s(n11595), .op(
        n5013) );
  mux2_1 U14147 ( .ip1(\cache_data[14][27] ), .ip2(n11642), .s(n11595), .op(
        n5012) );
  mux2_1 U14148 ( .ip1(\cache_data[14][28] ), .ip2(n11643), .s(n11595), .op(
        n5011) );
  mux2_1 U14149 ( .ip1(\cache_data[14][29] ), .ip2(n11644), .s(n11595), .op(
        n5010) );
  mux2_1 U14150 ( .ip1(\cache_data[14][30] ), .ip2(n11645), .s(n11595), .op(
        n5009) );
  mux2_1 U14151 ( .ip1(\cache_data[14][31] ), .ip2(n11647), .s(n11595), .op(
        n5008) );
  nor2_1 U14152 ( .ip1(n11606), .ip2(n11600), .op(n11596) );
  mux2_1 U14153 ( .ip1(\cache_data[14][32] ), .ip2(n11614), .s(n11596), .op(
        n5007) );
  mux2_1 U14154 ( .ip1(\cache_data[14][33] ), .ip2(n11615), .s(n11596), .op(
        n5006) );
  mux2_1 U14155 ( .ip1(\cache_data[14][34] ), .ip2(n11616), .s(n11596), .op(
        n5005) );
  mux2_1 U14156 ( .ip1(\cache_data[14][35] ), .ip2(n11617), .s(n11596), .op(
        n5004) );
  mux2_1 U14157 ( .ip1(\cache_data[14][36] ), .ip2(n11618), .s(n11596), .op(
        n5003) );
  mux2_1 U14158 ( .ip1(\cache_data[14][37] ), .ip2(n11619), .s(n11596), .op(
        n5002) );
  mux2_1 U14159 ( .ip1(\cache_data[14][38] ), .ip2(n11620), .s(n11596), .op(
        n5001) );
  mux2_1 U14160 ( .ip1(\cache_data[14][39] ), .ip2(n11621), .s(n11596), .op(
        n5000) );
  mux2_1 U14161 ( .ip1(\cache_data[14][40] ), .ip2(n11622), .s(n11596), .op(
        n4999) );
  mux2_1 U14162 ( .ip1(\cache_data[14][41] ), .ip2(n11623), .s(n11596), .op(
        n4998) );
  mux2_1 U14163 ( .ip1(\cache_data[14][42] ), .ip2(n11624), .s(n11596), .op(
        n4997) );
  mux2_1 U14164 ( .ip1(\cache_data[14][43] ), .ip2(n11625), .s(n11596), .op(
        n4996) );
  mux2_1 U14165 ( .ip1(\cache_data[14][44] ), .ip2(n11626), .s(n11596), .op(
        n4995) );
  mux2_1 U14166 ( .ip1(\cache_data[14][45] ), .ip2(n11627), .s(n11596), .op(
        n4994) );
  mux2_1 U14167 ( .ip1(\cache_data[14][46] ), .ip2(n11628), .s(n11596), .op(
        n4993) );
  mux2_1 U14168 ( .ip1(\cache_data[14][47] ), .ip2(n11629), .s(n11596), .op(
        n4992) );
  mux2_1 U14169 ( .ip1(\cache_data[14][48] ), .ip2(n11630), .s(n11596), .op(
        n4991) );
  mux2_1 U14170 ( .ip1(\cache_data[14][49] ), .ip2(n11631), .s(n11596), .op(
        n4990) );
  mux2_1 U14171 ( .ip1(\cache_data[14][50] ), .ip2(n11632), .s(n11596), .op(
        n4989) );
  buf_1 U14172 ( .ip(n11596), .op(n11597) );
  mux2_1 U14173 ( .ip1(\cache_data[14][51] ), .ip2(n11633), .s(n11597), .op(
        n4988) );
  mux2_1 U14174 ( .ip1(\cache_data[14][52] ), .ip2(n11634), .s(n11597), .op(
        n4987) );
  mux2_1 U14175 ( .ip1(\cache_data[14][53] ), .ip2(n11635), .s(n11597), .op(
        n4986) );
  mux2_1 U14176 ( .ip1(\cache_data[14][54] ), .ip2(n11636), .s(n11597), .op(
        n4985) );
  mux2_1 U14177 ( .ip1(\cache_data[14][55] ), .ip2(n11637), .s(n11597), .op(
        n4984) );
  mux2_1 U14178 ( .ip1(\cache_data[14][56] ), .ip2(n11638), .s(n11596), .op(
        n4983) );
  mux2_1 U14179 ( .ip1(\cache_data[14][57] ), .ip2(n11640), .s(n11596), .op(
        n4982) );
  mux2_1 U14180 ( .ip1(\cache_data[14][58] ), .ip2(n11641), .s(n11597), .op(
        n4981) );
  mux2_1 U14181 ( .ip1(\cache_data[14][59] ), .ip2(n11642), .s(n11597), .op(
        n4980) );
  mux2_1 U14182 ( .ip1(\cache_data[14][60] ), .ip2(n11643), .s(n11597), .op(
        n4979) );
  mux2_1 U14183 ( .ip1(\cache_data[14][61] ), .ip2(n11644), .s(n11597), .op(
        n4978) );
  mux2_1 U14184 ( .ip1(\cache_data[14][62] ), .ip2(n11645), .s(n11597), .op(
        n4977) );
  mux2_1 U14185 ( .ip1(\cache_data[14][63] ), .ip2(n11647), .s(n11597), .op(
        n4976) );
  nor2_1 U14186 ( .ip1(n11609), .ip2(n11600), .op(n11598) );
  mux2_1 U14187 ( .ip1(\cache_data[14][64] ), .ip2(n11614), .s(n11598), .op(
        n4975) );
  mux2_1 U14188 ( .ip1(\cache_data[14][65] ), .ip2(n11615), .s(n11598), .op(
        n4974) );
  mux2_1 U14189 ( .ip1(\cache_data[14][66] ), .ip2(n11616), .s(n11598), .op(
        n4973) );
  mux2_1 U14190 ( .ip1(\cache_data[14][67] ), .ip2(n11617), .s(n11598), .op(
        n4972) );
  mux2_1 U14191 ( .ip1(\cache_data[14][68] ), .ip2(n11618), .s(n11598), .op(
        n4971) );
  mux2_1 U14192 ( .ip1(\cache_data[14][69] ), .ip2(n11619), .s(n11598), .op(
        n4970) );
  mux2_1 U14193 ( .ip1(\cache_data[14][70] ), .ip2(n11620), .s(n11598), .op(
        n4969) );
  mux2_1 U14194 ( .ip1(\cache_data[14][71] ), .ip2(n11621), .s(n11598), .op(
        n4968) );
  mux2_1 U14195 ( .ip1(\cache_data[14][72] ), .ip2(n11622), .s(n11598), .op(
        n4967) );
  buf_1 U14196 ( .ip(n11598), .op(n11599) );
  mux2_1 U14197 ( .ip1(\cache_data[14][73] ), .ip2(n11623), .s(n11599), .op(
        n4966) );
  mux2_1 U14198 ( .ip1(\cache_data[14][74] ), .ip2(n11624), .s(n11599), .op(
        n4965) );
  mux2_1 U14199 ( .ip1(\cache_data[14][75] ), .ip2(n11625), .s(n11598), .op(
        n4964) );
  mux2_1 U14200 ( .ip1(\cache_data[14][76] ), .ip2(n11626), .s(n11598), .op(
        n4963) );
  mux2_1 U14201 ( .ip1(\cache_data[14][77] ), .ip2(n11627), .s(n11599), .op(
        n4962) );
  mux2_1 U14202 ( .ip1(\cache_data[14][78] ), .ip2(n11628), .s(n11598), .op(
        n4961) );
  mux2_1 U14203 ( .ip1(\cache_data[14][79] ), .ip2(n11629), .s(n11598), .op(
        n4960) );
  mux2_1 U14204 ( .ip1(\cache_data[14][80] ), .ip2(n11630), .s(n11598), .op(
        n4959) );
  mux2_1 U14205 ( .ip1(\cache_data[14][81] ), .ip2(n11631), .s(n11598), .op(
        n4958) );
  mux2_1 U14206 ( .ip1(\cache_data[14][82] ), .ip2(n11632), .s(n11598), .op(
        n4957) );
  mux2_1 U14207 ( .ip1(\cache_data[14][83] ), .ip2(n11633), .s(n11598), .op(
        n4956) );
  mux2_1 U14208 ( .ip1(\cache_data[14][84] ), .ip2(n11634), .s(n11598), .op(
        n4955) );
  mux2_1 U14209 ( .ip1(\cache_data[14][85] ), .ip2(n11635), .s(n11598), .op(
        n4954) );
  mux2_1 U14210 ( .ip1(\cache_data[14][86] ), .ip2(n11636), .s(n11598), .op(
        n4953) );
  mux2_1 U14211 ( .ip1(\cache_data[14][87] ), .ip2(n11637), .s(n11598), .op(
        n4952) );
  mux2_1 U14212 ( .ip1(\cache_data[14][88] ), .ip2(n11638), .s(n11599), .op(
        n4951) );
  mux2_1 U14213 ( .ip1(\cache_data[14][89] ), .ip2(n11640), .s(n11599), .op(
        n4950) );
  mux2_1 U14214 ( .ip1(\cache_data[14][90] ), .ip2(n11641), .s(n11599), .op(
        n4949) );
  mux2_1 U14215 ( .ip1(\cache_data[14][91] ), .ip2(n11642), .s(n11599), .op(
        n4948) );
  mux2_1 U14216 ( .ip1(\cache_data[14][92] ), .ip2(n11643), .s(n11599), .op(
        n4947) );
  mux2_1 U14217 ( .ip1(\cache_data[14][93] ), .ip2(n11644), .s(n11599), .op(
        n4946) );
  mux2_1 U14218 ( .ip1(\cache_data[14][94] ), .ip2(n11645), .s(n11599), .op(
        n4945) );
  mux2_1 U14219 ( .ip1(\cache_data[14][95] ), .ip2(n11647), .s(n11599), .op(
        n4944) );
  nor2_1 U14220 ( .ip1(n11613), .ip2(n11600), .op(n11601) );
  mux2_1 U14221 ( .ip1(\cache_data[14][96] ), .ip2(n11614), .s(n11601), .op(
        n4943) );
  mux2_1 U14222 ( .ip1(\cache_data[14][97] ), .ip2(n11615), .s(n11601), .op(
        n4942) );
  mux2_1 U14223 ( .ip1(\cache_data[14][98] ), .ip2(n11616), .s(n11601), .op(
        n4941) );
  mux2_1 U14224 ( .ip1(\cache_data[14][99] ), .ip2(n11617), .s(n11601), .op(
        n4940) );
  mux2_1 U14225 ( .ip1(\cache_data[14][100] ), .ip2(n11618), .s(n11601), .op(
        n4939) );
  mux2_1 U14226 ( .ip1(\cache_data[14][101] ), .ip2(n11619), .s(n11601), .op(
        n4938) );
  mux2_1 U14227 ( .ip1(\cache_data[14][102] ), .ip2(n11620), .s(n11601), .op(
        n4937) );
  mux2_1 U14228 ( .ip1(\cache_data[14][103] ), .ip2(n11621), .s(n11601), .op(
        n4936) );
  mux2_1 U14229 ( .ip1(\cache_data[14][104] ), .ip2(n11622), .s(n11601), .op(
        n4935) );
  buf_1 U14230 ( .ip(n11601), .op(n11602) );
  mux2_1 U14231 ( .ip1(\cache_data[14][105] ), .ip2(n11623), .s(n11602), .op(
        n4934) );
  mux2_1 U14232 ( .ip1(\cache_data[14][106] ), .ip2(n11624), .s(n11602), .op(
        n4933) );
  mux2_1 U14233 ( .ip1(\cache_data[14][107] ), .ip2(n11625), .s(n11601), .op(
        n4932) );
  mux2_1 U14234 ( .ip1(\cache_data[14][108] ), .ip2(n11626), .s(n11601), .op(
        n4931) );
  mux2_1 U14235 ( .ip1(\cache_data[14][109] ), .ip2(n11627), .s(n11602), .op(
        n4930) );
  mux2_1 U14236 ( .ip1(\cache_data[14][110] ), .ip2(n11628), .s(n11601), .op(
        n4929) );
  mux2_1 U14237 ( .ip1(\cache_data[14][111] ), .ip2(n11629), .s(n11601), .op(
        n4928) );
  mux2_1 U14238 ( .ip1(\cache_data[14][112] ), .ip2(n11630), .s(n11601), .op(
        n4927) );
  mux2_1 U14239 ( .ip1(\cache_data[14][113] ), .ip2(n11631), .s(n11601), .op(
        n4926) );
  mux2_1 U14240 ( .ip1(\cache_data[14][114] ), .ip2(n11632), .s(n11601), .op(
        n4925) );
  mux2_1 U14241 ( .ip1(\cache_data[14][115] ), .ip2(n11633), .s(n11601), .op(
        n4924) );
  mux2_1 U14242 ( .ip1(\cache_data[14][116] ), .ip2(n11634), .s(n11601), .op(
        n4923) );
  mux2_1 U14243 ( .ip1(\cache_data[14][117] ), .ip2(n11635), .s(n11601), .op(
        n4922) );
  mux2_1 U14244 ( .ip1(\cache_data[14][118] ), .ip2(n11636), .s(n11601), .op(
        n4921) );
  mux2_1 U14245 ( .ip1(\cache_data[14][119] ), .ip2(n11637), .s(n11601), .op(
        n4920) );
  mux2_1 U14246 ( .ip1(\cache_data[14][120] ), .ip2(n11638), .s(n11602), .op(
        n4919) );
  mux2_1 U14247 ( .ip1(\cache_data[14][121] ), .ip2(n11640), .s(n11602), .op(
        n4918) );
  mux2_1 U14248 ( .ip1(\cache_data[14][122] ), .ip2(n11641), .s(n11602), .op(
        n4917) );
  mux2_1 U14249 ( .ip1(\cache_data[14][123] ), .ip2(n11642), .s(n11602), .op(
        n4916) );
  mux2_1 U14250 ( .ip1(\cache_data[14][124] ), .ip2(n11643), .s(n11602), .op(
        n4915) );
  mux2_1 U14251 ( .ip1(\cache_data[14][125] ), .ip2(n11644), .s(n11602), .op(
        n4914) );
  mux2_1 U14252 ( .ip1(\cache_data[14][126] ), .ip2(n11645), .s(n11602), .op(
        n4913) );
  mux2_1 U14253 ( .ip1(\cache_data[14][127] ), .ip2(n11647), .s(n11602), .op(
        n4912) );
  nor2_1 U14254 ( .ip1(n11603), .ip2(n11612), .op(n11604) );
  mux2_1 U14255 ( .ip1(\cache_data[15][0] ), .ip2(n11614), .s(n11604), .op(
        n4911) );
  mux2_1 U14256 ( .ip1(\cache_data[15][1] ), .ip2(n11615), .s(n11604), .op(
        n4910) );
  mux2_1 U14257 ( .ip1(\cache_data[15][2] ), .ip2(n11616), .s(n11604), .op(
        n4909) );
  mux2_1 U14258 ( .ip1(\cache_data[15][3] ), .ip2(n11617), .s(n11604), .op(
        n4908) );
  mux2_1 U14259 ( .ip1(\cache_data[15][4] ), .ip2(n11618), .s(n11604), .op(
        n4907) );
  mux2_1 U14260 ( .ip1(\cache_data[15][5] ), .ip2(n11619), .s(n11604), .op(
        n4906) );
  mux2_1 U14261 ( .ip1(\cache_data[15][6] ), .ip2(n11620), .s(n11604), .op(
        n4905) );
  mux2_1 U14262 ( .ip1(\cache_data[15][7] ), .ip2(n11621), .s(n11604), .op(
        n4904) );
  mux2_1 U14263 ( .ip1(\cache_data[15][8] ), .ip2(n11622), .s(n11604), .op(
        n4903) );
  mux2_1 U14264 ( .ip1(\cache_data[15][9] ), .ip2(n11623), .s(n11604), .op(
        n4902) );
  mux2_1 U14265 ( .ip1(\cache_data[15][10] ), .ip2(n11624), .s(n11604), .op(
        n4901) );
  mux2_1 U14266 ( .ip1(\cache_data[15][11] ), .ip2(n11625), .s(n11604), .op(
        n4900) );
  mux2_1 U14267 ( .ip1(\cache_data[15][12] ), .ip2(n11626), .s(n11604), .op(
        n4899) );
  mux2_1 U14268 ( .ip1(\cache_data[15][13] ), .ip2(n11627), .s(n11604), .op(
        n4898) );
  mux2_1 U14269 ( .ip1(\cache_data[15][14] ), .ip2(n11628), .s(n11604), .op(
        n4897) );
  mux2_1 U14270 ( .ip1(\cache_data[15][15] ), .ip2(n11629), .s(n11604), .op(
        n4896) );
  mux2_1 U14271 ( .ip1(\cache_data[15][16] ), .ip2(n11630), .s(n11604), .op(
        n4895) );
  mux2_1 U14272 ( .ip1(\cache_data[15][17] ), .ip2(n11631), .s(n11604), .op(
        n4894) );
  mux2_1 U14273 ( .ip1(\cache_data[15][18] ), .ip2(n11632), .s(n11604), .op(
        n4893) );
  buf_1 U14274 ( .ip(n11604), .op(n11605) );
  mux2_1 U14275 ( .ip1(\cache_data[15][19] ), .ip2(n11633), .s(n11605), .op(
        n4892) );
  mux2_1 U14276 ( .ip1(\cache_data[15][20] ), .ip2(n11634), .s(n11605), .op(
        n4891) );
  mux2_1 U14277 ( .ip1(\cache_data[15][21] ), .ip2(n11635), .s(n11605), .op(
        n4890) );
  mux2_1 U14278 ( .ip1(\cache_data[15][22] ), .ip2(n11636), .s(n11605), .op(
        n4889) );
  mux2_1 U14279 ( .ip1(\cache_data[15][23] ), .ip2(n11637), .s(n11605), .op(
        n4888) );
  mux2_1 U14280 ( .ip1(\cache_data[15][24] ), .ip2(n11638), .s(n11604), .op(
        n4887) );
  mux2_1 U14281 ( .ip1(\cache_data[15][25] ), .ip2(n11640), .s(n11604), .op(
        n4886) );
  mux2_1 U14282 ( .ip1(\cache_data[15][26] ), .ip2(n11641), .s(n11605), .op(
        n4885) );
  mux2_1 U14283 ( .ip1(\cache_data[15][27] ), .ip2(n11642), .s(n11605), .op(
        n4884) );
  mux2_1 U14284 ( .ip1(\cache_data[15][28] ), .ip2(n11643), .s(n11605), .op(
        n4883) );
  mux2_1 U14285 ( .ip1(\cache_data[15][29] ), .ip2(n11644), .s(n11605), .op(
        n4882) );
  mux2_1 U14286 ( .ip1(\cache_data[15][30] ), .ip2(n11645), .s(n11605), .op(
        n4881) );
  mux2_1 U14287 ( .ip1(\cache_data[15][31] ), .ip2(n11647), .s(n11605), .op(
        n4880) );
  nor2_1 U14288 ( .ip1(n11606), .ip2(n11612), .op(n11607) );
  mux2_1 U14289 ( .ip1(\cache_data[15][32] ), .ip2(n11614), .s(n11607), .op(
        n4879) );
  mux2_1 U14290 ( .ip1(\cache_data[15][33] ), .ip2(n11615), .s(n11607), .op(
        n4878) );
  mux2_1 U14291 ( .ip1(\cache_data[15][34] ), .ip2(n11616), .s(n11607), .op(
        n4877) );
  mux2_1 U14292 ( .ip1(\cache_data[15][35] ), .ip2(n11617), .s(n11607), .op(
        n4876) );
  mux2_1 U14293 ( .ip1(\cache_data[15][36] ), .ip2(n11618), .s(n11607), .op(
        n4875) );
  mux2_1 U14294 ( .ip1(\cache_data[15][37] ), .ip2(n11619), .s(n11607), .op(
        n4874) );
  mux2_1 U14295 ( .ip1(\cache_data[15][38] ), .ip2(n11620), .s(n11607), .op(
        n4873) );
  mux2_1 U14296 ( .ip1(\cache_data[15][39] ), .ip2(n11621), .s(n11607), .op(
        n4872) );
  mux2_1 U14297 ( .ip1(\cache_data[15][40] ), .ip2(n11622), .s(n11607), .op(
        n4871) );
  mux2_1 U14298 ( .ip1(\cache_data[15][41] ), .ip2(n11623), .s(n11607), .op(
        n4870) );
  mux2_1 U14299 ( .ip1(\cache_data[15][42] ), .ip2(n11624), .s(n11607), .op(
        n4869) );
  mux2_1 U14300 ( .ip1(\cache_data[15][43] ), .ip2(n11625), .s(n11607), .op(
        n4868) );
  mux2_1 U14301 ( .ip1(\cache_data[15][44] ), .ip2(n11626), .s(n11607), .op(
        n4867) );
  mux2_1 U14302 ( .ip1(\cache_data[15][45] ), .ip2(n11627), .s(n11607), .op(
        n4866) );
  mux2_1 U14303 ( .ip1(\cache_data[15][46] ), .ip2(n11628), .s(n11607), .op(
        n4865) );
  mux2_1 U14304 ( .ip1(\cache_data[15][47] ), .ip2(n11629), .s(n11607), .op(
        n4864) );
  mux2_1 U14305 ( .ip1(\cache_data[15][48] ), .ip2(n11630), .s(n11607), .op(
        n4863) );
  mux2_1 U14306 ( .ip1(\cache_data[15][49] ), .ip2(n11631), .s(n11607), .op(
        n4862) );
  mux2_1 U14307 ( .ip1(\cache_data[15][50] ), .ip2(n11632), .s(n11607), .op(
        n4861) );
  buf_1 U14308 ( .ip(n11607), .op(n11608) );
  mux2_1 U14309 ( .ip1(\cache_data[15][51] ), .ip2(n11633), .s(n11608), .op(
        n4860) );
  mux2_1 U14310 ( .ip1(\cache_data[15][52] ), .ip2(n11634), .s(n11608), .op(
        n4859) );
  mux2_1 U14311 ( .ip1(\cache_data[15][53] ), .ip2(n11635), .s(n11608), .op(
        n4858) );
  mux2_1 U14312 ( .ip1(\cache_data[15][54] ), .ip2(n11636), .s(n11608), .op(
        n4857) );
  mux2_1 U14313 ( .ip1(\cache_data[15][55] ), .ip2(n11637), .s(n11608), .op(
        n4856) );
  mux2_1 U14314 ( .ip1(\cache_data[15][56] ), .ip2(n11638), .s(n11607), .op(
        n4855) );
  mux2_1 U14315 ( .ip1(\cache_data[15][57] ), .ip2(n11640), .s(n11607), .op(
        n4854) );
  mux2_1 U14316 ( .ip1(\cache_data[15][58] ), .ip2(n11641), .s(n11608), .op(
        n4853) );
  mux2_1 U14317 ( .ip1(\cache_data[15][59] ), .ip2(n11642), .s(n11608), .op(
        n4852) );
  mux2_1 U14318 ( .ip1(\cache_data[15][60] ), .ip2(n11643), .s(n11608), .op(
        n4851) );
  mux2_1 U14319 ( .ip1(\cache_data[15][61] ), .ip2(n11644), .s(n11608), .op(
        n4850) );
  mux2_1 U14320 ( .ip1(\cache_data[15][62] ), .ip2(n11645), .s(n11608), .op(
        n4849) );
  mux2_1 U14321 ( .ip1(\cache_data[15][63] ), .ip2(n11647), .s(n11608), .op(
        n4848) );
  nor2_1 U14322 ( .ip1(n11609), .ip2(n11612), .op(n11610) );
  mux2_1 U14323 ( .ip1(\cache_data[15][64] ), .ip2(n11614), .s(n11610), .op(
        n4847) );
  mux2_1 U14324 ( .ip1(\cache_data[15][65] ), .ip2(n11615), .s(n11610), .op(
        n4846) );
  mux2_1 U14325 ( .ip1(\cache_data[15][66] ), .ip2(n11616), .s(n11610), .op(
        n4845) );
  mux2_1 U14326 ( .ip1(\cache_data[15][67] ), .ip2(n11617), .s(n11610), .op(
        n4844) );
  mux2_1 U14327 ( .ip1(\cache_data[15][68] ), .ip2(n11618), .s(n11610), .op(
        n4843) );
  mux2_1 U14328 ( .ip1(\cache_data[15][69] ), .ip2(n11619), .s(n11610), .op(
        n4842) );
  mux2_1 U14329 ( .ip1(\cache_data[15][70] ), .ip2(n11620), .s(n11610), .op(
        n4841) );
  mux2_1 U14330 ( .ip1(\cache_data[15][71] ), .ip2(n11621), .s(n11610), .op(
        n4840) );
  mux2_1 U14331 ( .ip1(\cache_data[15][72] ), .ip2(n11622), .s(n11610), .op(
        n4839) );
  mux2_1 U14332 ( .ip1(\cache_data[15][73] ), .ip2(n11623), .s(n11610), .op(
        n4838) );
  mux2_1 U14333 ( .ip1(\cache_data[15][74] ), .ip2(n11624), .s(n11610), .op(
        n4837) );
  mux2_1 U14334 ( .ip1(\cache_data[15][75] ), .ip2(n11625), .s(n11610), .op(
        n4836) );
  mux2_1 U14335 ( .ip1(\cache_data[15][76] ), .ip2(n11626), .s(n11610), .op(
        n4835) );
  mux2_1 U14336 ( .ip1(\cache_data[15][77] ), .ip2(n11627), .s(n11610), .op(
        n4834) );
  mux2_1 U14337 ( .ip1(\cache_data[15][78] ), .ip2(n11628), .s(n11610), .op(
        n4833) );
  mux2_1 U14338 ( .ip1(\cache_data[15][79] ), .ip2(n11629), .s(n11610), .op(
        n4832) );
  mux2_1 U14339 ( .ip1(\cache_data[15][80] ), .ip2(n11630), .s(n11610), .op(
        n4831) );
  mux2_1 U14340 ( .ip1(\cache_data[15][81] ), .ip2(n11631), .s(n11610), .op(
        n4830) );
  mux2_1 U14341 ( .ip1(\cache_data[15][82] ), .ip2(n11632), .s(n11610), .op(
        n4829) );
  buf_1 U14342 ( .ip(n11610), .op(n11611) );
  mux2_1 U14343 ( .ip1(\cache_data[15][83] ), .ip2(n11633), .s(n11611), .op(
        n4828) );
  mux2_1 U14344 ( .ip1(\cache_data[15][84] ), .ip2(n11634), .s(n11611), .op(
        n4827) );
  mux2_1 U14345 ( .ip1(\cache_data[15][85] ), .ip2(n11635), .s(n11611), .op(
        n4826) );
  mux2_1 U14346 ( .ip1(\cache_data[15][86] ), .ip2(n11636), .s(n11611), .op(
        n4825) );
  mux2_1 U14347 ( .ip1(\cache_data[15][87] ), .ip2(n11637), .s(n11611), .op(
        n4824) );
  mux2_1 U14348 ( .ip1(\cache_data[15][88] ), .ip2(n11638), .s(n11610), .op(
        n4823) );
  mux2_1 U14349 ( .ip1(\cache_data[15][89] ), .ip2(n11640), .s(n11610), .op(
        n4822) );
  mux2_1 U14350 ( .ip1(\cache_data[15][90] ), .ip2(n11641), .s(n11611), .op(
        n4821) );
  mux2_1 U14351 ( .ip1(\cache_data[15][91] ), .ip2(n11642), .s(n11611), .op(
        n4820) );
  mux2_1 U14352 ( .ip1(\cache_data[15][92] ), .ip2(n11643), .s(n11611), .op(
        n4819) );
  mux2_1 U14353 ( .ip1(\cache_data[15][93] ), .ip2(n11644), .s(n11611), .op(
        n4818) );
  mux2_1 U14354 ( .ip1(\cache_data[15][94] ), .ip2(n11645), .s(n11611), .op(
        n4817) );
  mux2_1 U14355 ( .ip1(\cache_data[15][95] ), .ip2(n11647), .s(n11611), .op(
        n4816) );
  nor2_1 U14356 ( .ip1(n11613), .ip2(n11612), .op(n11639) );
  mux2_1 U14357 ( .ip1(\cache_data[15][96] ), .ip2(n11614), .s(n11639), .op(
        n4815) );
  mux2_1 U14358 ( .ip1(\cache_data[15][97] ), .ip2(n11615), .s(n11639), .op(
        n4814) );
  mux2_1 U14359 ( .ip1(\cache_data[15][98] ), .ip2(n11616), .s(n11639), .op(
        n4813) );
  mux2_1 U14360 ( .ip1(\cache_data[15][99] ), .ip2(n11617), .s(n11639), .op(
        n4812) );
  mux2_1 U14361 ( .ip1(\cache_data[15][100] ), .ip2(n11618), .s(n11639), .op(
        n4811) );
  mux2_1 U14362 ( .ip1(\cache_data[15][101] ), .ip2(n11619), .s(n11639), .op(
        n4810) );
  mux2_1 U14363 ( .ip1(\cache_data[15][102] ), .ip2(n11620), .s(n11639), .op(
        n4809) );
  mux2_1 U14364 ( .ip1(\cache_data[15][103] ), .ip2(n11621), .s(n11639), .op(
        n4808) );
  mux2_1 U14365 ( .ip1(\cache_data[15][104] ), .ip2(n11622), .s(n11639), .op(
        n4807) );
  mux2_1 U14366 ( .ip1(\cache_data[15][105] ), .ip2(n11623), .s(n11639), .op(
        n4806) );
  mux2_1 U14367 ( .ip1(\cache_data[15][106] ), .ip2(n11624), .s(n11639), .op(
        n4805) );
  mux2_1 U14368 ( .ip1(\cache_data[15][107] ), .ip2(n11625), .s(n11639), .op(
        n4804) );
  mux2_1 U14369 ( .ip1(\cache_data[15][108] ), .ip2(n11626), .s(n11639), .op(
        n4803) );
  mux2_1 U14370 ( .ip1(\cache_data[15][109] ), .ip2(n11627), .s(n11639), .op(
        n4802) );
  mux2_1 U14371 ( .ip1(\cache_data[15][110] ), .ip2(n11628), .s(n11639), .op(
        n4801) );
  mux2_1 U14372 ( .ip1(\cache_data[15][111] ), .ip2(n11629), .s(n11639), .op(
        n4800) );
  mux2_1 U14373 ( .ip1(\cache_data[15][112] ), .ip2(n11630), .s(n11639), .op(
        n4799) );
  mux2_1 U14374 ( .ip1(\cache_data[15][113] ), .ip2(n11631), .s(n11639), .op(
        n4798) );
  mux2_1 U14375 ( .ip1(\cache_data[15][114] ), .ip2(n11632), .s(n11639), .op(
        n4797) );
  buf_1 U14376 ( .ip(n11639), .op(n11646) );
  mux2_1 U14377 ( .ip1(\cache_data[15][115] ), .ip2(n11633), .s(n11646), .op(
        n4796) );
  mux2_1 U14378 ( .ip1(\cache_data[15][116] ), .ip2(n11634), .s(n11646), .op(
        n4795) );
  mux2_1 U14379 ( .ip1(\cache_data[15][117] ), .ip2(n11635), .s(n11646), .op(
        n4794) );
  mux2_1 U14380 ( .ip1(\cache_data[15][118] ), .ip2(n11636), .s(n11646), .op(
        n4793) );
  mux2_1 U14381 ( .ip1(\cache_data[15][119] ), .ip2(n11637), .s(n11646), .op(
        n4792) );
  mux2_1 U14382 ( .ip1(\cache_data[15][120] ), .ip2(n11638), .s(n11639), .op(
        n4791) );
  mux2_1 U14383 ( .ip1(\cache_data[15][121] ), .ip2(n11640), .s(n11639), .op(
        n4790) );
  mux2_1 U14384 ( .ip1(\cache_data[15][122] ), .ip2(n11641), .s(n11646), .op(
        n4789) );
  mux2_1 U14385 ( .ip1(\cache_data[15][123] ), .ip2(n11642), .s(n11646), .op(
        n4788) );
  mux2_1 U14386 ( .ip1(\cache_data[15][124] ), .ip2(n11643), .s(n11646), .op(
        n4787) );
  mux2_1 U14387 ( .ip1(\cache_data[15][125] ), .ip2(n11644), .s(n11646), .op(
        n4786) );
  mux2_1 U14388 ( .ip1(\cache_data[15][126] ), .ip2(n11645), .s(n11646), .op(
        n4785) );
  mux2_1 U14389 ( .ip1(\cache_data[15][127] ), .ip2(n11647), .s(n11646), .op(
        n4784) );
  nand2_1 U14390 ( .ip1(mem_data_cnt[2]), .ip2(n11658), .op(n11649) );
  nand2_1 U14391 ( .ip1(addr_mem[2]), .ip2(n12257), .op(n11648) );
  nand2_1 U14392 ( .ip1(n11649), .ip2(n11648), .op(n4781) );
  nand2_1 U14393 ( .ip1(mem_data_cnt[3]), .ip2(n11658), .op(n11651) );
  nand2_1 U14394 ( .ip1(addr_mem[3]), .ip2(n12257), .op(n11650) );
  nand2_1 U14395 ( .ip1(n11651), .ip2(n11650), .op(n4780) );
  nand2_1 U14396 ( .ip1(addr_resp[4]), .ip2(n11658), .op(n11653) );
  nand2_1 U14397 ( .ip1(addr_mem[4]), .ip2(n12257), .op(n11652) );
  nand2_1 U14398 ( .ip1(n11653), .ip2(n11652), .op(n4779) );
  nand2_1 U14399 ( .ip1(addr_resp[5]), .ip2(n11658), .op(n11655) );
  nand2_1 U14400 ( .ip1(addr_mem[5]), .ip2(n12257), .op(n11654) );
  nand2_1 U14401 ( .ip1(n11655), .ip2(n11654), .op(n4778) );
  nand2_1 U14402 ( .ip1(addr_resp[6]), .ip2(n11658), .op(n11657) );
  nand2_1 U14403 ( .ip1(addr_mem[6]), .ip2(n12257), .op(n11656) );
  nand2_1 U14404 ( .ip1(n11657), .ip2(n11656), .op(n4777) );
  nand2_1 U14405 ( .ip1(addr_resp[7]), .ip2(n11658), .op(n11660) );
  nand2_1 U14406 ( .ip1(addr_mem[7]), .ip2(n12257), .op(n11659) );
  nand2_1 U14407 ( .ip1(n11660), .ip2(n11659), .op(n4776) );
  nand2_1 U14408 ( .ip1(n11964), .ip2(\cache_tag[0][0] ), .op(n11664) );
  nand2_1 U14409 ( .ip1(n12170), .ip2(\cache_tag[11][0] ), .op(n11663) );
  nand2_1 U14410 ( .ip1(n12202), .ip2(\cache_tag[7][0] ), .op(n11662) );
  nand2_1 U14411 ( .ip1(n11965), .ip2(\cache_tag[15][0] ), .op(n11661) );
  nand4_1 U14412 ( .ip1(n11664), .ip2(n11663), .ip3(n11662), .ip4(n11661), 
        .op(n11680) );
  nand2_1 U14413 ( .ip1(n12234), .ip2(\cache_tag[8][0] ), .op(n11668) );
  nand2_1 U14414 ( .ip1(n11972), .ip2(\cache_tag[6][0] ), .op(n11667) );
  nand2_1 U14415 ( .ip1(n12242), .ip2(\cache_tag[13][0] ), .op(n11666) );
  nand2_1 U14416 ( .ip1(n11966), .ip2(\cache_tag[10][0] ), .op(n11665) );
  nand4_1 U14417 ( .ip1(n11668), .ip2(n11667), .ip3(n11666), .ip4(n11665), 
        .op(n11679) );
  nand2_1 U14418 ( .ip1(n12241), .ip2(\cache_tag[9][0] ), .op(n11672) );
  nand2_1 U14419 ( .ip1(n12030), .ip2(\cache_tag[12][0] ), .op(n11671) );
  nand2_1 U14420 ( .ip1(n11963), .ip2(\cache_tag[5][0] ), .op(n11670) );
  nand2_1 U14421 ( .ip1(n11973), .ip2(\cache_tag[2][0] ), .op(n11669) );
  nand4_1 U14422 ( .ip1(n11672), .ip2(n11671), .ip3(n11670), .ip4(n11669), 
        .op(n11678) );
  nand2_1 U14423 ( .ip1(n12164), .ip2(\cache_tag[4][0] ), .op(n11676) );
  nand2_1 U14424 ( .ip1(n11978), .ip2(\cache_tag[3][0] ), .op(n11675) );
  nand2_1 U14425 ( .ip1(n11688), .ip2(\cache_tag[14][0] ), .op(n11674) );
  nand2_1 U14426 ( .ip1(n11943), .ip2(\cache_tag[1][0] ), .op(n11673) );
  nand4_1 U14427 ( .ip1(n11676), .ip2(n11675), .ip3(n11674), .ip4(n11673), 
        .op(n11677) );
  nor4_1 U14428 ( .ip1(n11680), .ip2(n11679), .ip3(n11678), .ip4(n11677), .op(
        n11681) );
  nor2_1 U14429 ( .ip1(n11681), .ip2(n12252), .op(n11683) );
  and2_1 U14430 ( .ip1(n12254), .ip2(addr_resp[8]), .op(n11682) );
  ab_or_c_or_d U14431 ( .ip1(addr_mem[8]), .ip2(n12257), .ip3(n11683), .ip4(
        n11682), .op(n4775) );
  nand2_1 U14432 ( .ip1(n11978), .ip2(\cache_tag[3][1] ), .op(n11687) );
  nand2_1 U14433 ( .ip1(n11966), .ip2(\cache_tag[10][1] ), .op(n11686) );
  nand2_1 U14434 ( .ip1(n11963), .ip2(\cache_tag[5][1] ), .op(n11685) );
  nand2_1 U14435 ( .ip1(n12164), .ip2(\cache_tag[4][1] ), .op(n11684) );
  nand4_1 U14436 ( .ip1(n11687), .ip2(n11686), .ip3(n11685), .ip4(n11684), 
        .op(n11704) );
  nand2_1 U14437 ( .ip1(n11965), .ip2(\cache_tag[15][1] ), .op(n11692) );
  nand2_1 U14438 ( .ip1(n11688), .ip2(\cache_tag[14][1] ), .op(n11691) );
  nand2_1 U14439 ( .ip1(n12242), .ip2(\cache_tag[13][1] ), .op(n11690) );
  nand2_1 U14440 ( .ip1(n12170), .ip2(\cache_tag[11][1] ), .op(n11689) );
  nand4_1 U14441 ( .ip1(n11692), .ip2(n11691), .ip3(n11690), .ip4(n11689), 
        .op(n11703) );
  nand2_1 U14442 ( .ip1(n11979), .ip2(\cache_tag[1][1] ), .op(n11696) );
  nand2_1 U14443 ( .ip1(n12234), .ip2(\cache_tag[8][1] ), .op(n11695) );
  nand2_1 U14444 ( .ip1(n11972), .ip2(\cache_tag[6][1] ), .op(n11694) );
  nand2_1 U14445 ( .ip1(n12030), .ip2(\cache_tag[12][1] ), .op(n11693) );
  nand4_1 U14446 ( .ip1(n11696), .ip2(n11695), .ip3(n11694), .ip4(n11693), 
        .op(n11702) );
  nand2_1 U14447 ( .ip1(n11973), .ip2(\cache_tag[2][1] ), .op(n11700) );
  nand2_1 U14448 ( .ip1(n12241), .ip2(\cache_tag[9][1] ), .op(n11699) );
  nand2_1 U14449 ( .ip1(n12202), .ip2(\cache_tag[7][1] ), .op(n11698) );
  nand2_1 U14450 ( .ip1(n11964), .ip2(\cache_tag[0][1] ), .op(n11697) );
  nand4_1 U14451 ( .ip1(n11700), .ip2(n11699), .ip3(n11698), .ip4(n11697), 
        .op(n11701) );
  nor4_1 U14452 ( .ip1(n11704), .ip2(n11703), .ip3(n11702), .ip4(n11701), .op(
        n11705) );
  nor2_1 U14453 ( .ip1(n11705), .ip2(n12252), .op(n11707) );
  and2_1 U14454 ( .ip1(n12254), .ip2(addr_resp[9]), .op(n11706) );
  ab_or_c_or_d U14455 ( .ip1(addr_mem[9]), .ip2(n12257), .ip3(n11707), .ip4(
        n11706), .op(n4774) );
  nand2_1 U14456 ( .ip1(n11965), .ip2(\cache_tag[15][2] ), .op(n11711) );
  nand2_1 U14457 ( .ip1(n11971), .ip2(\cache_tag[14][2] ), .op(n11710) );
  nand2_1 U14458 ( .ip1(n11927), .ip2(\cache_tag[11][2] ), .op(n11709) );
  nand2_1 U14459 ( .ip1(n12164), .ip2(\cache_tag[4][2] ), .op(n11708) );
  nand4_1 U14460 ( .ip1(n11711), .ip2(n11710), .ip3(n11709), .ip4(n11708), 
        .op(n11727) );
  nand2_1 U14461 ( .ip1(n11973), .ip2(\cache_tag[2][2] ), .op(n11715) );
  nand2_1 U14462 ( .ip1(n11979), .ip2(\cache_tag[1][2] ), .op(n11714) );
  nand2_1 U14463 ( .ip1(n11963), .ip2(\cache_tag[5][2] ), .op(n11713) );
  nand2_1 U14464 ( .ip1(n11972), .ip2(\cache_tag[6][2] ), .op(n11712) );
  nand4_1 U14465 ( .ip1(n11715), .ip2(n11714), .ip3(n11713), .ip4(n11712), 
        .op(n11726) );
  nand2_1 U14466 ( .ip1(n12234), .ip2(\cache_tag[8][2] ), .op(n11719) );
  nand2_1 U14467 ( .ip1(n11966), .ip2(\cache_tag[10][2] ), .op(n11718) );
  nand2_1 U14468 ( .ip1(n11978), .ip2(\cache_tag[3][2] ), .op(n11717) );
  nand2_1 U14469 ( .ip1(n12242), .ip2(\cache_tag[13][2] ), .op(n11716) );
  nand4_1 U14470 ( .ip1(n11719), .ip2(n11718), .ip3(n11717), .ip4(n11716), 
        .op(n11725) );
  nand2_1 U14471 ( .ip1(n12030), .ip2(\cache_tag[12][2] ), .op(n11723) );
  nand2_1 U14472 ( .ip1(n11964), .ip2(\cache_tag[0][2] ), .op(n11722) );
  nand2_1 U14473 ( .ip1(n12152), .ip2(\cache_tag[9][2] ), .op(n11721) );
  nand2_1 U14474 ( .ip1(n12202), .ip2(\cache_tag[7][2] ), .op(n11720) );
  nand4_1 U14475 ( .ip1(n11723), .ip2(n11722), .ip3(n11721), .ip4(n11720), 
        .op(n11724) );
  nor4_1 U14476 ( .ip1(n11727), .ip2(n11726), .ip3(n11725), .ip4(n11724), .op(
        n11728) );
  nor2_1 U14477 ( .ip1(n11728), .ip2(n12252), .op(n11730) );
  and2_1 U14478 ( .ip1(n12254), .ip2(addr_resp[10]), .op(n11729) );
  ab_or_c_or_d U14479 ( .ip1(addr_mem[10]), .ip2(n12257), .ip3(n11730), .ip4(
        n11729), .op(n4773) );
  nand2_1 U14480 ( .ip1(n12227), .ip2(\cache_tag[12][3] ), .op(n11734) );
  nand2_1 U14481 ( .ip1(n11971), .ip2(\cache_tag[14][3] ), .op(n11733) );
  nand2_1 U14482 ( .ip1(n11964), .ip2(\cache_tag[0][3] ), .op(n11732) );
  nand2_1 U14483 ( .ip1(n12241), .ip2(\cache_tag[9][3] ), .op(n11731) );
  nand4_1 U14484 ( .ip1(n11734), .ip2(n11733), .ip3(n11732), .ip4(n11731), 
        .op(n11750) );
  nand2_1 U14485 ( .ip1(n11943), .ip2(\cache_tag[1][3] ), .op(n11738) );
  nand2_1 U14486 ( .ip1(n11978), .ip2(\cache_tag[3][3] ), .op(n11737) );
  nand2_1 U14487 ( .ip1(n12170), .ip2(\cache_tag[11][3] ), .op(n11736) );
  nand2_1 U14488 ( .ip1(n11966), .ip2(\cache_tag[10][3] ), .op(n11735) );
  nand4_1 U14489 ( .ip1(n11738), .ip2(n11737), .ip3(n11736), .ip4(n11735), 
        .op(n11749) );
  nand2_1 U14490 ( .ip1(n11963), .ip2(\cache_tag[5][3] ), .op(n11742) );
  nand2_1 U14491 ( .ip1(n11965), .ip2(\cache_tag[15][3] ), .op(n11741) );
  nand2_1 U14492 ( .ip1(n11973), .ip2(\cache_tag[2][3] ), .op(n11740) );
  nand2_1 U14493 ( .ip1(n12165), .ip2(\cache_tag[13][3] ), .op(n11739) );
  nand4_1 U14494 ( .ip1(n11742), .ip2(n11741), .ip3(n11740), .ip4(n11739), 
        .op(n11748) );
  nand2_1 U14495 ( .ip1(n12191), .ip2(\cache_tag[8][3] ), .op(n11746) );
  nand2_1 U14496 ( .ip1(n12143), .ip2(\cache_tag[7][3] ), .op(n11745) );
  nand2_1 U14497 ( .ip1(n11972), .ip2(\cache_tag[6][3] ), .op(n11744) );
  nand2_1 U14498 ( .ip1(n12164), .ip2(\cache_tag[4][3] ), .op(n11743) );
  nand4_1 U14499 ( .ip1(n11746), .ip2(n11745), .ip3(n11744), .ip4(n11743), 
        .op(n11747) );
  nor4_1 U14500 ( .ip1(n11750), .ip2(n11749), .ip3(n11748), .ip4(n11747), .op(
        n11751) );
  nor2_1 U14501 ( .ip1(n11751), .ip2(n12252), .op(n11753) );
  and2_1 U14502 ( .ip1(n12254), .ip2(addr_resp[11]), .op(n11752) );
  ab_or_c_or_d U14503 ( .ip1(addr_mem[11]), .ip2(n12257), .ip3(n11753), .ip4(
        n11752), .op(n4772) );
  nand2_1 U14504 ( .ip1(n11978), .ip2(\cache_tag[3][4] ), .op(n11757) );
  nand2_1 U14505 ( .ip1(n11971), .ip2(\cache_tag[14][4] ), .op(n11756) );
  nand2_1 U14506 ( .ip1(n11972), .ip2(\cache_tag[6][4] ), .op(n11755) );
  nand2_1 U14507 ( .ip1(n11966), .ip2(\cache_tag[10][4] ), .op(n11754) );
  nand4_1 U14508 ( .ip1(n11757), .ip2(n11756), .ip3(n11755), .ip4(n11754), 
        .op(n11773) );
  nand2_1 U14509 ( .ip1(n11973), .ip2(\cache_tag[2][4] ), .op(n11761) );
  nand2_1 U14510 ( .ip1(n11963), .ip2(\cache_tag[5][4] ), .op(n11760) );
  nand2_1 U14511 ( .ip1(n11943), .ip2(\cache_tag[1][4] ), .op(n11759) );
  nand2_1 U14512 ( .ip1(n11964), .ip2(\cache_tag[0][4] ), .op(n11758) );
  nand4_1 U14513 ( .ip1(n11761), .ip2(n11760), .ip3(n11759), .ip4(n11758), 
        .op(n11772) );
  nand2_1 U14514 ( .ip1(n12143), .ip2(\cache_tag[7][4] ), .op(n11765) );
  nand2_1 U14515 ( .ip1(n11965), .ip2(\cache_tag[15][4] ), .op(n11764) );
  nand2_1 U14516 ( .ip1(n12164), .ip2(\cache_tag[4][4] ), .op(n11763) );
  nand2_1 U14517 ( .ip1(n12242), .ip2(\cache_tag[13][4] ), .op(n11762) );
  nand4_1 U14518 ( .ip1(n11765), .ip2(n11764), .ip3(n11763), .ip4(n11762), 
        .op(n11771) );
  nand2_1 U14519 ( .ip1(n12030), .ip2(\cache_tag[12][4] ), .op(n11769) );
  nand2_1 U14520 ( .ip1(n12152), .ip2(\cache_tag[9][4] ), .op(n11768) );
  nand2_1 U14521 ( .ip1(n12191), .ip2(\cache_tag[8][4] ), .op(n11767) );
  nand2_1 U14522 ( .ip1(n12170), .ip2(\cache_tag[11][4] ), .op(n11766) );
  nand4_1 U14523 ( .ip1(n11769), .ip2(n11768), .ip3(n11767), .ip4(n11766), 
        .op(n11770) );
  nor4_1 U14524 ( .ip1(n11773), .ip2(n11772), .ip3(n11771), .ip4(n11770), .op(
        n11774) );
  nor2_1 U14525 ( .ip1(n11774), .ip2(n12252), .op(n11776) );
  and2_1 U14526 ( .ip1(n12254), .ip2(addr_resp[12]), .op(n11775) );
  ab_or_c_or_d U14527 ( .ip1(addr_mem[12]), .ip2(n12257), .ip3(n11776), .ip4(
        n11775), .op(n4771) );
  nand2_1 U14528 ( .ip1(n12152), .ip2(\cache_tag[9][5] ), .op(n11780) );
  nand2_1 U14529 ( .ip1(n11979), .ip2(\cache_tag[1][5] ), .op(n11779) );
  nand2_1 U14530 ( .ip1(n12165), .ip2(\cache_tag[13][5] ), .op(n11778) );
  nand2_1 U14531 ( .ip1(n12202), .ip2(\cache_tag[7][5] ), .op(n11777) );
  nand4_1 U14532 ( .ip1(n11780), .ip2(n11779), .ip3(n11778), .ip4(n11777), 
        .op(n11796) );
  nand2_1 U14533 ( .ip1(n11971), .ip2(\cache_tag[14][5] ), .op(n11784) );
  nand2_1 U14534 ( .ip1(n11973), .ip2(\cache_tag[2][5] ), .op(n11783) );
  nand2_1 U14535 ( .ip1(n11964), .ip2(\cache_tag[0][5] ), .op(n11782) );
  nand2_1 U14536 ( .ip1(n12164), .ip2(\cache_tag[4][5] ), .op(n11781) );
  nand4_1 U14537 ( .ip1(n11784), .ip2(n11783), .ip3(n11782), .ip4(n11781), 
        .op(n11795) );
  nand2_1 U14538 ( .ip1(n12030), .ip2(\cache_tag[12][5] ), .op(n11788) );
  nand2_1 U14539 ( .ip1(n11963), .ip2(\cache_tag[5][5] ), .op(n11787) );
  nand2_1 U14540 ( .ip1(n12191), .ip2(\cache_tag[8][5] ), .op(n11786) );
  nand2_1 U14541 ( .ip1(n11978), .ip2(\cache_tag[3][5] ), .op(n11785) );
  nand4_1 U14542 ( .ip1(n11788), .ip2(n11787), .ip3(n11786), .ip4(n11785), 
        .op(n11794) );
  nand2_1 U14543 ( .ip1(n11972), .ip2(\cache_tag[6][5] ), .op(n11792) );
  nand2_1 U14544 ( .ip1(n11965), .ip2(\cache_tag[15][5] ), .op(n11791) );
  nand2_1 U14545 ( .ip1(n11927), .ip2(\cache_tag[11][5] ), .op(n11790) );
  nand2_1 U14546 ( .ip1(n11966), .ip2(\cache_tag[10][5] ), .op(n11789) );
  nand4_1 U14547 ( .ip1(n11792), .ip2(n11791), .ip3(n11790), .ip4(n11789), 
        .op(n11793) );
  nor4_1 U14548 ( .ip1(n11796), .ip2(n11795), .ip3(n11794), .ip4(n11793), .op(
        n11797) );
  nor2_1 U14549 ( .ip1(n11797), .ip2(n12252), .op(n11799) );
  and2_1 U14550 ( .ip1(n12254), .ip2(addr_resp[13]), .op(n11798) );
  ab_or_c_or_d U14551 ( .ip1(addr_mem[13]), .ip2(n12257), .ip3(n11799), .ip4(
        n11798), .op(n4770) );
  nand2_1 U14552 ( .ip1(n11966), .ip2(\cache_tag[10][6] ), .op(n11803) );
  nand2_1 U14553 ( .ip1(n11963), .ip2(\cache_tag[5][6] ), .op(n11802) );
  nand2_1 U14554 ( .ip1(n11978), .ip2(\cache_tag[3][6] ), .op(n11801) );
  nand2_1 U14555 ( .ip1(n12234), .ip2(\cache_tag[8][6] ), .op(n11800) );
  nand4_1 U14556 ( .ip1(n11803), .ip2(n11802), .ip3(n11801), .ip4(n11800), 
        .op(n11819) );
  nand2_1 U14557 ( .ip1(n11964), .ip2(\cache_tag[0][6] ), .op(n11807) );
  nand2_1 U14558 ( .ip1(n11972), .ip2(\cache_tag[6][6] ), .op(n11806) );
  nand2_1 U14559 ( .ip1(n11973), .ip2(\cache_tag[2][6] ), .op(n11805) );
  nand2_1 U14560 ( .ip1(n12242), .ip2(\cache_tag[13][6] ), .op(n11804) );
  nand4_1 U14561 ( .ip1(n11807), .ip2(n11806), .ip3(n11805), .ip4(n11804), 
        .op(n11818) );
  nand2_1 U14562 ( .ip1(n12170), .ip2(\cache_tag[11][6] ), .op(n11811) );
  nand2_1 U14563 ( .ip1(n11971), .ip2(\cache_tag[14][6] ), .op(n11810) );
  nand2_1 U14564 ( .ip1(n12241), .ip2(\cache_tag[9][6] ), .op(n11809) );
  nand2_1 U14565 ( .ip1(n12030), .ip2(\cache_tag[12][6] ), .op(n11808) );
  nand4_1 U14566 ( .ip1(n11811), .ip2(n11810), .ip3(n11809), .ip4(n11808), 
        .op(n11817) );
  nand2_1 U14567 ( .ip1(n11965), .ip2(\cache_tag[15][6] ), .op(n11815) );
  nand2_1 U14568 ( .ip1(n12164), .ip2(\cache_tag[4][6] ), .op(n11814) );
  nand2_1 U14569 ( .ip1(n11979), .ip2(\cache_tag[1][6] ), .op(n11813) );
  nand2_1 U14570 ( .ip1(n12143), .ip2(\cache_tag[7][6] ), .op(n11812) );
  nand4_1 U14571 ( .ip1(n11815), .ip2(n11814), .ip3(n11813), .ip4(n11812), 
        .op(n11816) );
  nor4_1 U14572 ( .ip1(n11819), .ip2(n11818), .ip3(n11817), .ip4(n11816), .op(
        n11820) );
  nor2_1 U14573 ( .ip1(n11820), .ip2(n12252), .op(n11822) );
  and2_1 U14574 ( .ip1(n12254), .ip2(addr_resp[14]), .op(n11821) );
  ab_or_c_or_d U14575 ( .ip1(addr_mem[14]), .ip2(n12257), .ip3(n11822), .ip4(
        n11821), .op(n4769) );
  nand2_1 U14576 ( .ip1(n12243), .ip2(\cache_tag[4][7] ), .op(n11826) );
  nand2_1 U14577 ( .ip1(n12152), .ip2(\cache_tag[9][7] ), .op(n11825) );
  nand2_1 U14578 ( .ip1(n11943), .ip2(\cache_tag[1][7] ), .op(n11824) );
  nand2_1 U14579 ( .ip1(n11973), .ip2(\cache_tag[2][7] ), .op(n11823) );
  nand4_1 U14580 ( .ip1(n11826), .ip2(n11825), .ip3(n11824), .ip4(n11823), 
        .op(n11842) );
  nand2_1 U14581 ( .ip1(n11965), .ip2(\cache_tag[15][7] ), .op(n11830) );
  nand2_1 U14582 ( .ip1(n11966), .ip2(\cache_tag[10][7] ), .op(n11829) );
  nand2_1 U14583 ( .ip1(n11978), .ip2(\cache_tag[3][7] ), .op(n11828) );
  nand2_1 U14584 ( .ip1(n12170), .ip2(\cache_tag[11][7] ), .op(n11827) );
  nand4_1 U14585 ( .ip1(n11830), .ip2(n11829), .ip3(n11828), .ip4(n11827), 
        .op(n11841) );
  nand2_1 U14586 ( .ip1(n12234), .ip2(\cache_tag[8][7] ), .op(n11834) );
  nand2_1 U14587 ( .ip1(n11964), .ip2(\cache_tag[0][7] ), .op(n11833) );
  nand2_1 U14588 ( .ip1(n11972), .ip2(\cache_tag[6][7] ), .op(n11832) );
  nand2_1 U14589 ( .ip1(n12242), .ip2(\cache_tag[13][7] ), .op(n11831) );
  nand4_1 U14590 ( .ip1(n11834), .ip2(n11833), .ip3(n11832), .ip4(n11831), 
        .op(n11840) );
  nand2_1 U14591 ( .ip1(n11971), .ip2(\cache_tag[14][7] ), .op(n11838) );
  nand2_1 U14592 ( .ip1(n11963), .ip2(\cache_tag[5][7] ), .op(n11837) );
  nand2_1 U14593 ( .ip1(n12030), .ip2(\cache_tag[12][7] ), .op(n11836) );
  nand2_1 U14594 ( .ip1(n12143), .ip2(\cache_tag[7][7] ), .op(n11835) );
  nand4_1 U14595 ( .ip1(n11838), .ip2(n11837), .ip3(n11836), .ip4(n11835), 
        .op(n11839) );
  nor4_1 U14596 ( .ip1(n11842), .ip2(n11841), .ip3(n11840), .ip4(n11839), .op(
        n11843) );
  nor2_1 U14597 ( .ip1(n11843), .ip2(n12252), .op(n11845) );
  and2_1 U14598 ( .ip1(n12254), .ip2(addr_resp[15]), .op(n11844) );
  ab_or_c_or_d U14599 ( .ip1(addr_mem[15]), .ip2(n12257), .ip3(n11845), .ip4(
        n11844), .op(n4768) );
  nand2_1 U14600 ( .ip1(n12152), .ip2(\cache_tag[9][8] ), .op(n11849) );
  nand2_1 U14601 ( .ip1(n11927), .ip2(\cache_tag[11][8] ), .op(n11848) );
  nand2_1 U14602 ( .ip1(n12202), .ip2(\cache_tag[7][8] ), .op(n11847) );
  nand2_1 U14603 ( .ip1(n11971), .ip2(\cache_tag[14][8] ), .op(n11846) );
  nand4_1 U14604 ( .ip1(n11849), .ip2(n11848), .ip3(n11847), .ip4(n11846), 
        .op(n11865) );
  nand2_1 U14605 ( .ip1(n11972), .ip2(\cache_tag[6][8] ), .op(n11853) );
  nand2_1 U14606 ( .ip1(n11979), .ip2(\cache_tag[1][8] ), .op(n11852) );
  nand2_1 U14607 ( .ip1(n11965), .ip2(\cache_tag[15][8] ), .op(n11851) );
  nand2_1 U14608 ( .ip1(n11973), .ip2(\cache_tag[2][8] ), .op(n11850) );
  nand4_1 U14609 ( .ip1(n11853), .ip2(n11852), .ip3(n11851), .ip4(n11850), 
        .op(n11864) );
  nand2_1 U14610 ( .ip1(n11966), .ip2(\cache_tag[10][8] ), .op(n11857) );
  nand2_1 U14611 ( .ip1(n12164), .ip2(\cache_tag[4][8] ), .op(n11856) );
  nand2_1 U14612 ( .ip1(n11964), .ip2(\cache_tag[0][8] ), .op(n11855) );
  nand2_1 U14613 ( .ip1(n11963), .ip2(\cache_tag[5][8] ), .op(n11854) );
  nand4_1 U14614 ( .ip1(n11857), .ip2(n11856), .ip3(n11855), .ip4(n11854), 
        .op(n11863) );
  nand2_1 U14615 ( .ip1(n12030), .ip2(\cache_tag[12][8] ), .op(n11861) );
  nand2_1 U14616 ( .ip1(n12234), .ip2(\cache_tag[8][8] ), .op(n11860) );
  nand2_1 U14617 ( .ip1(n12165), .ip2(\cache_tag[13][8] ), .op(n11859) );
  nand2_1 U14618 ( .ip1(n11978), .ip2(\cache_tag[3][8] ), .op(n11858) );
  nand4_1 U14619 ( .ip1(n11861), .ip2(n11860), .ip3(n11859), .ip4(n11858), 
        .op(n11862) );
  nor4_1 U14620 ( .ip1(n11865), .ip2(n11864), .ip3(n11863), .ip4(n11862), .op(
        n11866) );
  nor2_1 U14621 ( .ip1(n11866), .ip2(n12252), .op(n11868) );
  and2_1 U14622 ( .ip1(n12254), .ip2(addr_resp[16]), .op(n11867) );
  ab_or_c_or_d U14623 ( .ip1(addr_mem[16]), .ip2(n12257), .ip3(n11868), .ip4(
        n11867), .op(n4767) );
  nand2_1 U14624 ( .ip1(n12241), .ip2(\cache_tag[9][9] ), .op(n11872) );
  nand2_1 U14625 ( .ip1(n12143), .ip2(\cache_tag[7][9] ), .op(n11871) );
  nand2_1 U14626 ( .ip1(n11963), .ip2(\cache_tag[5][9] ), .op(n11870) );
  nand2_1 U14627 ( .ip1(n11972), .ip2(\cache_tag[6][9] ), .op(n11869) );
  nand4_1 U14628 ( .ip1(n11872), .ip2(n11871), .ip3(n11870), .ip4(n11869), 
        .op(n11888) );
  nand2_1 U14629 ( .ip1(n12243), .ip2(\cache_tag[4][9] ), .op(n11876) );
  nand2_1 U14630 ( .ip1(n12165), .ip2(\cache_tag[13][9] ), .op(n11875) );
  nand2_1 U14631 ( .ip1(n12170), .ip2(\cache_tag[11][9] ), .op(n11874) );
  nand2_1 U14632 ( .ip1(n11965), .ip2(\cache_tag[15][9] ), .op(n11873) );
  nand4_1 U14633 ( .ip1(n11876), .ip2(n11875), .ip3(n11874), .ip4(n11873), 
        .op(n11887) );
  nand2_1 U14634 ( .ip1(n11966), .ip2(\cache_tag[10][9] ), .op(n11880) );
  nand2_1 U14635 ( .ip1(n11971), .ip2(\cache_tag[14][9] ), .op(n11879) );
  nand2_1 U14636 ( .ip1(n11973), .ip2(\cache_tag[2][9] ), .op(n11878) );
  nand2_1 U14637 ( .ip1(n11964), .ip2(\cache_tag[0][9] ), .op(n11877) );
  nand4_1 U14638 ( .ip1(n11880), .ip2(n11879), .ip3(n11878), .ip4(n11877), 
        .op(n11886) );
  nand2_1 U14639 ( .ip1(n12227), .ip2(\cache_tag[12][9] ), .op(n11884) );
  nand2_1 U14640 ( .ip1(n12234), .ip2(\cache_tag[8][9] ), .op(n11883) );
  nand2_1 U14641 ( .ip1(n11943), .ip2(\cache_tag[1][9] ), .op(n11882) );
  nand2_1 U14642 ( .ip1(n11978), .ip2(\cache_tag[3][9] ), .op(n11881) );
  nand4_1 U14643 ( .ip1(n11884), .ip2(n11883), .ip3(n11882), .ip4(n11881), 
        .op(n11885) );
  nor4_1 U14644 ( .ip1(n11888), .ip2(n11887), .ip3(n11886), .ip4(n11885), .op(
        n11889) );
  nor2_1 U14645 ( .ip1(n11889), .ip2(n12252), .op(n11891) );
  and2_1 U14646 ( .ip1(n12254), .ip2(addr_resp[17]), .op(n11890) );
  ab_or_c_or_d U14647 ( .ip1(addr_mem[17]), .ip2(n12257), .ip3(n11891), .ip4(
        n11890), .op(n4766) );
  nand2_1 U14648 ( .ip1(n11966), .ip2(\cache_tag[10][10] ), .op(n11895) );
  nand2_1 U14649 ( .ip1(n12152), .ip2(\cache_tag[9][10] ), .op(n11894) );
  nand2_1 U14650 ( .ip1(n11972), .ip2(\cache_tag[6][10] ), .op(n11893) );
  nand2_1 U14651 ( .ip1(n11943), .ip2(\cache_tag[1][10] ), .op(n11892) );
  nand4_1 U14652 ( .ip1(n11895), .ip2(n11894), .ip3(n11893), .ip4(n11892), 
        .op(n11911) );
  nand2_1 U14653 ( .ip1(n12170), .ip2(\cache_tag[11][10] ), .op(n11899) );
  nand2_1 U14654 ( .ip1(n11978), .ip2(\cache_tag[3][10] ), .op(n11898) );
  nand2_1 U14655 ( .ip1(n11963), .ip2(\cache_tag[5][10] ), .op(n11897) );
  nand2_1 U14656 ( .ip1(n12143), .ip2(\cache_tag[7][10] ), .op(n11896) );
  nand4_1 U14657 ( .ip1(n11899), .ip2(n11898), .ip3(n11897), .ip4(n11896), 
        .op(n11910) );
  nand2_1 U14658 ( .ip1(n11965), .ip2(\cache_tag[15][10] ), .op(n11903) );
  nand2_1 U14659 ( .ip1(n12164), .ip2(\cache_tag[4][10] ), .op(n11902) );
  nand2_1 U14660 ( .ip1(n11973), .ip2(\cache_tag[2][10] ), .op(n11901) );
  nand2_1 U14661 ( .ip1(n12234), .ip2(\cache_tag[8][10] ), .op(n11900) );
  nand4_1 U14662 ( .ip1(n11903), .ip2(n11902), .ip3(n11901), .ip4(n11900), 
        .op(n11909) );
  nand2_1 U14663 ( .ip1(n11964), .ip2(\cache_tag[0][10] ), .op(n11907) );
  nand2_1 U14664 ( .ip1(n12030), .ip2(\cache_tag[12][10] ), .op(n11906) );
  nand2_1 U14665 ( .ip1(n12242), .ip2(\cache_tag[13][10] ), .op(n11905) );
  nand2_1 U14666 ( .ip1(n11971), .ip2(\cache_tag[14][10] ), .op(n11904) );
  nand4_1 U14667 ( .ip1(n11907), .ip2(n11906), .ip3(n11905), .ip4(n11904), 
        .op(n11908) );
  nor4_1 U14668 ( .ip1(n11911), .ip2(n11910), .ip3(n11909), .ip4(n11908), .op(
        n11912) );
  nor2_1 U14669 ( .ip1(n11912), .ip2(n12252), .op(n11914) );
  and2_1 U14670 ( .ip1(n12254), .ip2(addr_resp[18]), .op(n11913) );
  ab_or_c_or_d U14671 ( .ip1(addr_mem[18]), .ip2(n12257), .ip3(n11914), .ip4(
        n11913), .op(n4765) );
  nand2_1 U14672 ( .ip1(n11978), .ip2(\cache_tag[3][11] ), .op(n11918) );
  nand2_1 U14673 ( .ip1(n12152), .ip2(\cache_tag[9][11] ), .op(n11917) );
  nand2_1 U14674 ( .ip1(n11971), .ip2(\cache_tag[14][11] ), .op(n11916) );
  nand2_1 U14675 ( .ip1(n12234), .ip2(\cache_tag[8][11] ), .op(n11915) );
  nand4_1 U14676 ( .ip1(n11918), .ip2(n11917), .ip3(n11916), .ip4(n11915), 
        .op(n11935) );
  nand2_1 U14677 ( .ip1(n12227), .ip2(\cache_tag[12][11] ), .op(n11922) );
  nand2_1 U14678 ( .ip1(n11973), .ip2(\cache_tag[2][11] ), .op(n11921) );
  nand2_1 U14679 ( .ip1(n12202), .ip2(\cache_tag[7][11] ), .op(n11920) );
  nand2_1 U14680 ( .ip1(n11966), .ip2(\cache_tag[10][11] ), .op(n11919) );
  nand4_1 U14681 ( .ip1(n11922), .ip2(n11921), .ip3(n11920), .ip4(n11919), 
        .op(n11934) );
  nand2_1 U14682 ( .ip1(n12165), .ip2(\cache_tag[13][11] ), .op(n11926) );
  nand2_1 U14683 ( .ip1(n12243), .ip2(\cache_tag[4][11] ), .op(n11925) );
  nand2_1 U14684 ( .ip1(n11979), .ip2(\cache_tag[1][11] ), .op(n11924) );
  nand2_1 U14685 ( .ip1(n11964), .ip2(\cache_tag[0][11] ), .op(n11923) );
  nand4_1 U14686 ( .ip1(n11926), .ip2(n11925), .ip3(n11924), .ip4(n11923), 
        .op(n11933) );
  nand2_1 U14687 ( .ip1(n11963), .ip2(\cache_tag[5][11] ), .op(n11931) );
  nand2_1 U14688 ( .ip1(n11927), .ip2(\cache_tag[11][11] ), .op(n11930) );
  nand2_1 U14689 ( .ip1(n11972), .ip2(\cache_tag[6][11] ), .op(n11929) );
  nand2_1 U14690 ( .ip1(n11965), .ip2(\cache_tag[15][11] ), .op(n11928) );
  nand4_1 U14691 ( .ip1(n11931), .ip2(n11930), .ip3(n11929), .ip4(n11928), 
        .op(n11932) );
  nor4_1 U14692 ( .ip1(n11935), .ip2(n11934), .ip3(n11933), .ip4(n11932), .op(
        n11936) );
  nor2_1 U14693 ( .ip1(n11936), .ip2(n12252), .op(n11938) );
  and2_1 U14694 ( .ip1(n12254), .ip2(addr_resp[19]), .op(n11937) );
  ab_or_c_or_d U14695 ( .ip1(addr_mem[19]), .ip2(n12257), .ip3(n11938), .ip4(
        n11937), .op(n4764) );
  nand2_1 U14696 ( .ip1(n12164), .ip2(\cache_tag[4][12] ), .op(n11942) );
  nand2_1 U14697 ( .ip1(n12030), .ip2(\cache_tag[12][12] ), .op(n11941) );
  nand2_1 U14698 ( .ip1(n12170), .ip2(\cache_tag[11][12] ), .op(n11940) );
  nand2_1 U14699 ( .ip1(n11966), .ip2(\cache_tag[10][12] ), .op(n11939) );
  nand4_1 U14700 ( .ip1(n11942), .ip2(n11941), .ip3(n11940), .ip4(n11939), 
        .op(n11959) );
  nand2_1 U14701 ( .ip1(n11963), .ip2(\cache_tag[5][12] ), .op(n11947) );
  nand2_1 U14702 ( .ip1(n11965), .ip2(\cache_tag[15][12] ), .op(n11946) );
  nand2_1 U14703 ( .ip1(n11943), .ip2(\cache_tag[1][12] ), .op(n11945) );
  nand2_1 U14704 ( .ip1(n12143), .ip2(\cache_tag[7][12] ), .op(n11944) );
  nand4_1 U14705 ( .ip1(n11947), .ip2(n11946), .ip3(n11945), .ip4(n11944), 
        .op(n11958) );
  nand2_1 U14706 ( .ip1(n12242), .ip2(\cache_tag[13][12] ), .op(n11951) );
  nand2_1 U14707 ( .ip1(n12241), .ip2(\cache_tag[9][12] ), .op(n11950) );
  nand2_1 U14708 ( .ip1(n11971), .ip2(\cache_tag[14][12] ), .op(n11949) );
  nand2_1 U14709 ( .ip1(n12191), .ip2(\cache_tag[8][12] ), .op(n11948) );
  nand4_1 U14710 ( .ip1(n11951), .ip2(n11950), .ip3(n11949), .ip4(n11948), 
        .op(n11957) );
  nand2_1 U14711 ( .ip1(n11964), .ip2(\cache_tag[0][12] ), .op(n11955) );
  nand2_1 U14712 ( .ip1(n11973), .ip2(\cache_tag[2][12] ), .op(n11954) );
  nand2_1 U14713 ( .ip1(n11972), .ip2(\cache_tag[6][12] ), .op(n11953) );
  nand2_1 U14714 ( .ip1(n11978), .ip2(\cache_tag[3][12] ), .op(n11952) );
  nand4_1 U14715 ( .ip1(n11955), .ip2(n11954), .ip3(n11953), .ip4(n11952), 
        .op(n11956) );
  nor4_1 U14716 ( .ip1(n11959), .ip2(n11958), .ip3(n11957), .ip4(n11956), .op(
        n11960) );
  nor2_1 U14717 ( .ip1(n11960), .ip2(n12252), .op(n11962) );
  and2_1 U14718 ( .ip1(n12254), .ip2(addr_resp[20]), .op(n11961) );
  ab_or_c_or_d U14719 ( .ip1(addr_mem[20]), .ip2(n12257), .ip3(n11962), .ip4(
        n11961), .op(n4763) );
  nand2_1 U14720 ( .ip1(n11963), .ip2(\cache_tag[5][13] ), .op(n11970) );
  nand2_1 U14721 ( .ip1(n11964), .ip2(\cache_tag[0][13] ), .op(n11969) );
  nand2_1 U14722 ( .ip1(n11965), .ip2(\cache_tag[15][13] ), .op(n11968) );
  nand2_1 U14723 ( .ip1(n11966), .ip2(\cache_tag[10][13] ), .op(n11967) );
  nand4_1 U14724 ( .ip1(n11970), .ip2(n11969), .ip3(n11968), .ip4(n11967), 
        .op(n11991) );
  nand2_1 U14725 ( .ip1(n12164), .ip2(\cache_tag[4][13] ), .op(n11977) );
  nand2_1 U14726 ( .ip1(n11971), .ip2(\cache_tag[14][13] ), .op(n11976) );
  nand2_1 U14727 ( .ip1(n11972), .ip2(\cache_tag[6][13] ), .op(n11975) );
  nand2_1 U14728 ( .ip1(n11973), .ip2(\cache_tag[2][13] ), .op(n11974) );
  nand4_1 U14729 ( .ip1(n11977), .ip2(n11976), .ip3(n11975), .ip4(n11974), 
        .op(n11990) );
  nand2_1 U14730 ( .ip1(n11978), .ip2(\cache_tag[3][13] ), .op(n11983) );
  nand2_1 U14731 ( .ip1(n12234), .ip2(\cache_tag[8][13] ), .op(n11982) );
  nand2_1 U14732 ( .ip1(n11979), .ip2(\cache_tag[1][13] ), .op(n11981) );
  nand2_1 U14733 ( .ip1(n12242), .ip2(\cache_tag[13][13] ), .op(n11980) );
  nand4_1 U14734 ( .ip1(n11983), .ip2(n11982), .ip3(n11981), .ip4(n11980), 
        .op(n11989) );
  nand2_1 U14735 ( .ip1(n12143), .ip2(\cache_tag[7][13] ), .op(n11987) );
  nand2_1 U14736 ( .ip1(n12170), .ip2(\cache_tag[11][13] ), .op(n11986) );
  nand2_1 U14737 ( .ip1(n12227), .ip2(\cache_tag[12][13] ), .op(n11985) );
  nand2_1 U14738 ( .ip1(n12152), .ip2(\cache_tag[9][13] ), .op(n11984) );
  nand4_1 U14739 ( .ip1(n11987), .ip2(n11986), .ip3(n11985), .ip4(n11984), 
        .op(n11988) );
  nor4_1 U14740 ( .ip1(n11991), .ip2(n11990), .ip3(n11989), .ip4(n11988), .op(
        n11992) );
  nor2_1 U14741 ( .ip1(n11992), .ip2(n12252), .op(n11994) );
  and2_1 U14742 ( .ip1(n12254), .ip2(addr_resp[21]), .op(n11993) );
  ab_or_c_or_d U14743 ( .ip1(addr_mem[21]), .ip2(n12257), .ip3(n11994), .ip4(
        n11993), .op(n4762) );
  nand2_1 U14744 ( .ip1(n12220), .ip2(\cache_tag[14][14] ), .op(n11998) );
  nand2_1 U14745 ( .ip1(n12219), .ip2(\cache_tag[3][14] ), .op(n11997) );
  nand2_1 U14746 ( .ip1(n12221), .ip2(\cache_tag[15][14] ), .op(n11996) );
  nand2_1 U14747 ( .ip1(n11979), .ip2(\cache_tag[1][14] ), .op(n11995) );
  nand4_1 U14748 ( .ip1(n11998), .ip2(n11997), .ip3(n11996), .ip4(n11995), 
        .op(n12014) );
  nand2_1 U14749 ( .ip1(n12121), .ip2(\cache_tag[8][14] ), .op(n12002) );
  nand2_1 U14750 ( .ip1(n12143), .ip2(\cache_tag[7][14] ), .op(n12001) );
  nand2_1 U14751 ( .ip1(n12096), .ip2(\cache_tag[11][14] ), .op(n12000) );
  nand2_1 U14752 ( .ip1(n12196), .ip2(\cache_tag[10][14] ), .op(n11999) );
  nand4_1 U14753 ( .ip1(n12002), .ip2(n12001), .ip3(n12000), .ip4(n11999), 
        .op(n12013) );
  nand2_1 U14754 ( .ip1(n12201), .ip2(\cache_tag[4][14] ), .op(n12006) );
  nand2_1 U14755 ( .ip1(n12030), .ip2(\cache_tag[12][14] ), .op(n12005) );
  nand2_1 U14756 ( .ip1(n12228), .ip2(\cache_tag[2][14] ), .op(n12004) );
  nand2_1 U14757 ( .ip1(n12233), .ip2(\cache_tag[0][14] ), .op(n12003) );
  nand4_1 U14758 ( .ip1(n12006), .ip2(n12005), .ip3(n12004), .ip4(n12003), 
        .op(n12012) );
  nand2_1 U14759 ( .ip1(n12142), .ip2(\cache_tag[13][14] ), .op(n12010) );
  nand2_1 U14760 ( .ip1(n10305), .ip2(\cache_tag[6][14] ), .op(n12009) );
  nand2_1 U14761 ( .ip1(n12241), .ip2(\cache_tag[9][14] ), .op(n12008) );
  nand2_1 U14762 ( .ip1(n12240), .ip2(\cache_tag[5][14] ), .op(n12007) );
  nand4_1 U14763 ( .ip1(n12010), .ip2(n12009), .ip3(n12008), .ip4(n12007), 
        .op(n12011) );
  nor4_1 U14764 ( .ip1(n12014), .ip2(n12013), .ip3(n12012), .ip4(n12011), .op(
        n12015) );
  nor2_1 U14765 ( .ip1(n12015), .ip2(n12252), .op(n12017) );
  and2_1 U14766 ( .ip1(n12254), .ip2(addr_resp[22]), .op(n12016) );
  ab_or_c_or_d U14767 ( .ip1(addr_mem[22]), .ip2(n12257), .ip3(n12017), .ip4(
        n12016), .op(n4761) );
  nand2_1 U14768 ( .ip1(n12142), .ip2(\cache_tag[13][15] ), .op(n12021) );
  nand2_1 U14769 ( .ip1(n12202), .ip2(\cache_tag[7][15] ), .op(n12020) );
  nand2_1 U14770 ( .ip1(n12096), .ip2(\cache_tag[11][15] ), .op(n12019) );
  nand2_1 U14771 ( .ip1(n12228), .ip2(\cache_tag[2][15] ), .op(n12018) );
  nand4_1 U14772 ( .ip1(n12021), .ip2(n12020), .ip3(n12019), .ip4(n12018), 
        .op(n12038) );
  nand2_1 U14773 ( .ip1(n12240), .ip2(\cache_tag[5][15] ), .op(n12025) );
  nand2_1 U14774 ( .ip1(n12243), .ip2(\cache_tag[4][15] ), .op(n12024) );
  nand2_1 U14775 ( .ip1(n12234), .ip2(\cache_tag[8][15] ), .op(n12023) );
  nand2_1 U14776 ( .ip1(n12233), .ip2(\cache_tag[0][15] ), .op(n12022) );
  nand4_1 U14777 ( .ip1(n12025), .ip2(n12024), .ip3(n12023), .ip4(n12022), 
        .op(n12037) );
  nand2_1 U14778 ( .ip1(n12126), .ip2(\cache_tag[9][15] ), .op(n12029) );
  nand2_1 U14779 ( .ip1(n12179), .ip2(\cache_tag[6][15] ), .op(n12028) );
  nand2_1 U14780 ( .ip1(n12196), .ip2(\cache_tag[10][15] ), .op(n12027) );
  nand2_1 U14781 ( .ip1(n12221), .ip2(\cache_tag[15][15] ), .op(n12026) );
  nand4_1 U14782 ( .ip1(n12029), .ip2(n12028), .ip3(n12027), .ip4(n12026), 
        .op(n12036) );
  nand2_1 U14783 ( .ip1(n12219), .ip2(\cache_tag[3][15] ), .op(n12034) );
  nand2_1 U14784 ( .ip1(n12220), .ip2(\cache_tag[14][15] ), .op(n12033) );
  nand2_1 U14785 ( .ip1(n12030), .ip2(\cache_tag[12][15] ), .op(n12032) );
  nand2_1 U14786 ( .ip1(n11943), .ip2(\cache_tag[1][15] ), .op(n12031) );
  nand4_1 U14787 ( .ip1(n12034), .ip2(n12033), .ip3(n12032), .ip4(n12031), 
        .op(n12035) );
  nor4_1 U14788 ( .ip1(n12038), .ip2(n12037), .ip3(n12036), .ip4(n12035), .op(
        n12039) );
  nor2_1 U14789 ( .ip1(n12039), .ip2(n12252), .op(n12041) );
  and2_1 U14790 ( .ip1(n12254), .ip2(addr_resp[23]), .op(n12040) );
  ab_or_c_or_d U14791 ( .ip1(addr_mem[23]), .ip2(n12257), .ip3(n12041), .ip4(
        n12040), .op(n4760) );
  nand2_1 U14792 ( .ip1(n12152), .ip2(\cache_tag[9][16] ), .op(n12045) );
  nand2_1 U14793 ( .ip1(n12219), .ip2(\cache_tag[3][16] ), .op(n12044) );
  nand2_1 U14794 ( .ip1(n11943), .ip2(\cache_tag[1][16] ), .op(n12043) );
  nand2_1 U14795 ( .ip1(n12191), .ip2(\cache_tag[8][16] ), .op(n12042) );
  nand4_1 U14796 ( .ip1(n12045), .ip2(n12044), .ip3(n12043), .ip4(n12042), 
        .op(n12061) );
  nand2_1 U14797 ( .ip1(n12221), .ip2(\cache_tag[15][16] ), .op(n12049) );
  nand2_1 U14798 ( .ip1(n12235), .ip2(\cache_tag[10][16] ), .op(n12048) );
  nand2_1 U14799 ( .ip1(n12233), .ip2(\cache_tag[0][16] ), .op(n12047) );
  nand2_1 U14800 ( .ip1(n12165), .ip2(\cache_tag[13][16] ), .op(n12046) );
  nand4_1 U14801 ( .ip1(n12049), .ip2(n12048), .ip3(n12047), .ip4(n12046), 
        .op(n12060) );
  nand2_1 U14802 ( .ip1(n10305), .ip2(\cache_tag[6][16] ), .op(n12053) );
  nand2_1 U14803 ( .ip1(n12096), .ip2(\cache_tag[11][16] ), .op(n12052) );
  nand2_1 U14804 ( .ip1(n12240), .ip2(\cache_tag[5][16] ), .op(n12051) );
  nand2_1 U14805 ( .ip1(n12243), .ip2(\cache_tag[4][16] ), .op(n12050) );
  nand4_1 U14806 ( .ip1(n12053), .ip2(n12052), .ip3(n12051), .ip4(n12050), 
        .op(n12059) );
  nand2_1 U14807 ( .ip1(n9560), .ip2(\cache_tag[12][16] ), .op(n12057) );
  nand2_1 U14808 ( .ip1(n12228), .ip2(\cache_tag[2][16] ), .op(n12056) );
  nand2_1 U14809 ( .ip1(n12202), .ip2(\cache_tag[7][16] ), .op(n12055) );
  nand2_1 U14810 ( .ip1(n12220), .ip2(\cache_tag[14][16] ), .op(n12054) );
  nand4_1 U14811 ( .ip1(n12057), .ip2(n12056), .ip3(n12055), .ip4(n12054), 
        .op(n12058) );
  nor4_1 U14812 ( .ip1(n12061), .ip2(n12060), .ip3(n12059), .ip4(n12058), .op(
        n12062) );
  nor2_1 U14813 ( .ip1(n12062), .ip2(n12252), .op(n12064) );
  and2_1 U14814 ( .ip1(n12254), .ip2(addr_resp[24]), .op(n12063) );
  ab_or_c_or_d U14815 ( .ip1(addr_mem[24]), .ip2(n12257), .ip3(n12064), .ip4(
        n12063), .op(n4759) );
  nand2_1 U14816 ( .ip1(n12220), .ip2(\cache_tag[14][17] ), .op(n12068) );
  nand2_1 U14817 ( .ip1(n12243), .ip2(\cache_tag[4][17] ), .op(n12067) );
  nand2_1 U14818 ( .ip1(n12165), .ip2(\cache_tag[13][17] ), .op(n12066) );
  nand2_1 U14819 ( .ip1(n12240), .ip2(\cache_tag[5][17] ), .op(n12065) );
  nand4_1 U14820 ( .ip1(n12068), .ip2(n12067), .ip3(n12066), .ip4(n12065), 
        .op(n12084) );
  nand2_1 U14821 ( .ip1(n12226), .ip2(\cache_tag[7][17] ), .op(n12072) );
  nand2_1 U14822 ( .ip1(n12241), .ip2(\cache_tag[9][17] ), .op(n12071) );
  nand2_1 U14823 ( .ip1(n12219), .ip2(\cache_tag[3][17] ), .op(n12070) );
  nand2_1 U14824 ( .ip1(n12235), .ip2(\cache_tag[10][17] ), .op(n12069) );
  nand4_1 U14825 ( .ip1(n12072), .ip2(n12071), .ip3(n12070), .ip4(n12069), 
        .op(n12083) );
  nand2_1 U14826 ( .ip1(n12228), .ip2(\cache_tag[2][17] ), .op(n12076) );
  nand2_1 U14827 ( .ip1(n9669), .ip2(\cache_tag[11][17] ), .op(n12075) );
  nand2_1 U14828 ( .ip1(n12233), .ip2(\cache_tag[0][17] ), .op(n12074) );
  nand2_1 U14829 ( .ip1(n12120), .ip2(\cache_tag[1][17] ), .op(n12073) );
  nand4_1 U14830 ( .ip1(n12076), .ip2(n12075), .ip3(n12074), .ip4(n12073), 
        .op(n12082) );
  nand2_1 U14831 ( .ip1(n12221), .ip2(\cache_tag[15][17] ), .op(n12080) );
  nand2_1 U14832 ( .ip1(n9560), .ip2(\cache_tag[12][17] ), .op(n12079) );
  nand2_1 U14833 ( .ip1(n12179), .ip2(\cache_tag[6][17] ), .op(n12078) );
  nand2_1 U14834 ( .ip1(n12191), .ip2(\cache_tag[8][17] ), .op(n12077) );
  nand4_1 U14835 ( .ip1(n12080), .ip2(n12079), .ip3(n12078), .ip4(n12077), 
        .op(n12081) );
  nor4_1 U14836 ( .ip1(n12084), .ip2(n12083), .ip3(n12082), .ip4(n12081), .op(
        n12085) );
  nor2_1 U14837 ( .ip1(n12085), .ip2(n12252), .op(n12087) );
  and2_1 U14838 ( .ip1(n12254), .ip2(addr_resp[25]), .op(n12086) );
  ab_or_c_or_d U14839 ( .ip1(addr_mem[25]), .ip2(n12257), .ip3(n12087), .ip4(
        n12086), .op(n4758) );
  nand2_1 U14840 ( .ip1(n12219), .ip2(\cache_tag[3][18] ), .op(n12091) );
  nand2_1 U14841 ( .ip1(n12240), .ip2(\cache_tag[5][18] ), .op(n12090) );
  nand2_1 U14842 ( .ip1(n9560), .ip2(\cache_tag[12][18] ), .op(n12089) );
  nand2_1 U14843 ( .ip1(n12191), .ip2(\cache_tag[8][18] ), .op(n12088) );
  nand4_1 U14844 ( .ip1(n12091), .ip2(n12090), .ip3(n12089), .ip4(n12088), 
        .op(n12108) );
  nand2_1 U14845 ( .ip1(n12233), .ip2(\cache_tag[0][18] ), .op(n12095) );
  nand2_1 U14846 ( .ip1(n12152), .ip2(\cache_tag[9][18] ), .op(n12094) );
  nand2_1 U14847 ( .ip1(n12235), .ip2(\cache_tag[10][18] ), .op(n12093) );
  nand2_1 U14848 ( .ip1(n11943), .ip2(\cache_tag[1][18] ), .op(n12092) );
  nand4_1 U14849 ( .ip1(n12095), .ip2(n12094), .ip3(n12093), .ip4(n12092), 
        .op(n12107) );
  nand2_1 U14850 ( .ip1(n12221), .ip2(\cache_tag[15][18] ), .op(n12100) );
  nand2_1 U14851 ( .ip1(n12096), .ip2(\cache_tag[11][18] ), .op(n12099) );
  nand2_1 U14852 ( .ip1(n12179), .ip2(\cache_tag[6][18] ), .op(n12098) );
  nand2_1 U14853 ( .ip1(n12228), .ip2(\cache_tag[2][18] ), .op(n12097) );
  nand4_1 U14854 ( .ip1(n12100), .ip2(n12099), .ip3(n12098), .ip4(n12097), 
        .op(n12106) );
  nand2_1 U14855 ( .ip1(n12164), .ip2(\cache_tag[4][18] ), .op(n12104) );
  nand2_1 U14856 ( .ip1(n12220), .ip2(\cache_tag[14][18] ), .op(n12103) );
  nand2_1 U14857 ( .ip1(n12202), .ip2(\cache_tag[7][18] ), .op(n12102) );
  nand2_1 U14858 ( .ip1(n12165), .ip2(\cache_tag[13][18] ), .op(n12101) );
  nand4_1 U14859 ( .ip1(n12104), .ip2(n12103), .ip3(n12102), .ip4(n12101), 
        .op(n12105) );
  nor4_1 U14860 ( .ip1(n12108), .ip2(n12107), .ip3(n12106), .ip4(n12105), .op(
        n12109) );
  nor2_1 U14861 ( .ip1(n12109), .ip2(n12252), .op(n12111) );
  and2_1 U14862 ( .ip1(n12254), .ip2(addr_resp[26]), .op(n12110) );
  ab_or_c_or_d U14863 ( .ip1(addr_mem[26]), .ip2(n12257), .ip3(n12111), .ip4(
        n12110), .op(n4757) );
  nand2_1 U14864 ( .ip1(n12233), .ip2(\cache_tag[0][19] ), .op(n12115) );
  nand2_1 U14865 ( .ip1(n12196), .ip2(\cache_tag[10][19] ), .op(n12114) );
  nand2_1 U14866 ( .ip1(n12170), .ip2(\cache_tag[11][19] ), .op(n12113) );
  nand2_1 U14867 ( .ip1(n12219), .ip2(\cache_tag[3][19] ), .op(n12112) );
  nand4_1 U14868 ( .ip1(n12115), .ip2(n12114), .ip3(n12113), .ip4(n12112), 
        .op(n12134) );
  nand2_1 U14869 ( .ip1(n12142), .ip2(\cache_tag[13][19] ), .op(n12119) );
  nand2_1 U14870 ( .ip1(n12179), .ip2(\cache_tag[6][19] ), .op(n12118) );
  nand2_1 U14871 ( .ip1(n12227), .ip2(\cache_tag[12][19] ), .op(n12117) );
  nand2_1 U14872 ( .ip1(n12240), .ip2(\cache_tag[5][19] ), .op(n12116) );
  nand4_1 U14873 ( .ip1(n12119), .ip2(n12118), .ip3(n12117), .ip4(n12116), 
        .op(n12133) );
  nand2_1 U14874 ( .ip1(n12221), .ip2(\cache_tag[15][19] ), .op(n12125) );
  nand2_1 U14875 ( .ip1(n12120), .ip2(\cache_tag[1][19] ), .op(n12124) );
  nand2_1 U14876 ( .ip1(n12121), .ip2(\cache_tag[8][19] ), .op(n12123) );
  nand2_1 U14877 ( .ip1(n12228), .ip2(\cache_tag[2][19] ), .op(n12122) );
  nand4_1 U14878 ( .ip1(n12125), .ip2(n12124), .ip3(n12123), .ip4(n12122), 
        .op(n12132) );
  nand2_1 U14879 ( .ip1(n12126), .ip2(\cache_tag[9][19] ), .op(n12130) );
  nand2_1 U14880 ( .ip1(n12220), .ip2(\cache_tag[14][19] ), .op(n12129) );
  nand2_1 U14881 ( .ip1(n12243), .ip2(\cache_tag[4][19] ), .op(n12128) );
  nand2_1 U14882 ( .ip1(n12202), .ip2(\cache_tag[7][19] ), .op(n12127) );
  nand4_1 U14883 ( .ip1(n12130), .ip2(n12129), .ip3(n12128), .ip4(n12127), 
        .op(n12131) );
  nor4_1 U14884 ( .ip1(n12134), .ip2(n12133), .ip3(n12132), .ip4(n12131), .op(
        n12135) );
  nor2_1 U14885 ( .ip1(n12135), .ip2(n12252), .op(n12137) );
  and2_1 U14886 ( .ip1(n12254), .ip2(addr_resp[27]), .op(n12136) );
  ab_or_c_or_d U14887 ( .ip1(addr_mem[27]), .ip2(n12257), .ip3(n12137), .ip4(
        n12136), .op(n4756) );
  nand2_1 U14888 ( .ip1(n12164), .ip2(\cache_tag[4][20] ), .op(n12141) );
  nand2_1 U14889 ( .ip1(n12221), .ip2(\cache_tag[15][20] ), .op(n12140) );
  nand2_1 U14890 ( .ip1(n11979), .ip2(\cache_tag[1][20] ), .op(n12139) );
  nand2_1 U14891 ( .ip1(n9669), .ip2(\cache_tag[11][20] ), .op(n12138) );
  nand4_1 U14892 ( .ip1(n12141), .ip2(n12140), .ip3(n12139), .ip4(n12138), 
        .op(n12160) );
  nand2_1 U14893 ( .ip1(n12142), .ip2(\cache_tag[13][20] ), .op(n12147) );
  nand2_1 U14894 ( .ip1(n12143), .ip2(\cache_tag[7][20] ), .op(n12146) );
  nand2_1 U14895 ( .ip1(n12235), .ip2(\cache_tag[10][20] ), .op(n12145) );
  nand2_1 U14896 ( .ip1(n12233), .ip2(\cache_tag[0][20] ), .op(n12144) );
  nand4_1 U14897 ( .ip1(n12147), .ip2(n12146), .ip3(n12145), .ip4(n12144), 
        .op(n12159) );
  nand2_1 U14898 ( .ip1(n12219), .ip2(\cache_tag[3][20] ), .op(n12151) );
  nand2_1 U14899 ( .ip1(n12234), .ip2(\cache_tag[8][20] ), .op(n12150) );
  nand2_1 U14900 ( .ip1(n12220), .ip2(\cache_tag[14][20] ), .op(n12149) );
  nand2_1 U14901 ( .ip1(n12179), .ip2(\cache_tag[6][20] ), .op(n12148) );
  nand4_1 U14902 ( .ip1(n12151), .ip2(n12150), .ip3(n12149), .ip4(n12148), 
        .op(n12158) );
  nand2_1 U14903 ( .ip1(n12207), .ip2(\cache_tag[12][20] ), .op(n12156) );
  nand2_1 U14904 ( .ip1(n12240), .ip2(\cache_tag[5][20] ), .op(n12155) );
  nand2_1 U14905 ( .ip1(n12152), .ip2(\cache_tag[9][20] ), .op(n12154) );
  nand2_1 U14906 ( .ip1(n12228), .ip2(\cache_tag[2][20] ), .op(n12153) );
  nand4_1 U14907 ( .ip1(n12156), .ip2(n12155), .ip3(n12154), .ip4(n12153), 
        .op(n12157) );
  nor4_1 U14908 ( .ip1(n12160), .ip2(n12159), .ip3(n12158), .ip4(n12157), .op(
        n12161) );
  nor2_1 U14909 ( .ip1(n12161), .ip2(n12252), .op(n12163) );
  and2_1 U14910 ( .ip1(n12254), .ip2(addr_resp[28]), .op(n12162) );
  ab_or_c_or_d U14911 ( .ip1(addr_mem[28]), .ip2(n12257), .ip3(n12163), .ip4(
        n12162), .op(n4755) );
  nand2_1 U14912 ( .ip1(n12164), .ip2(\cache_tag[4][21] ), .op(n12169) );
  nand2_1 U14913 ( .ip1(n12220), .ip2(\cache_tag[14][21] ), .op(n12168) );
  nand2_1 U14914 ( .ip1(n12191), .ip2(\cache_tag[8][21] ), .op(n12167) );
  nand2_1 U14915 ( .ip1(n12165), .ip2(\cache_tag[13][21] ), .op(n12166) );
  nand4_1 U14916 ( .ip1(n12169), .ip2(n12168), .ip3(n12167), .ip4(n12166), 
        .op(n12187) );
  nand2_1 U14917 ( .ip1(n12219), .ip2(\cache_tag[3][21] ), .op(n12174) );
  nand2_1 U14918 ( .ip1(n12170), .ip2(\cache_tag[11][21] ), .op(n12173) );
  nand2_1 U14919 ( .ip1(n12241), .ip2(\cache_tag[9][21] ), .op(n12172) );
  nand2_1 U14920 ( .ip1(n12240), .ip2(\cache_tag[5][21] ), .op(n12171) );
  nand4_1 U14921 ( .ip1(n12174), .ip2(n12173), .ip3(n12172), .ip4(n12171), 
        .op(n12186) );
  nand2_1 U14922 ( .ip1(n12226), .ip2(\cache_tag[7][21] ), .op(n12178) );
  nand2_1 U14923 ( .ip1(n12221), .ip2(\cache_tag[15][21] ), .op(n12177) );
  nand2_1 U14924 ( .ip1(n11979), .ip2(\cache_tag[1][21] ), .op(n12176) );
  nand2_1 U14925 ( .ip1(n12228), .ip2(\cache_tag[2][21] ), .op(n12175) );
  nand4_1 U14926 ( .ip1(n12178), .ip2(n12177), .ip3(n12176), .ip4(n12175), 
        .op(n12185) );
  nand2_1 U14927 ( .ip1(n9560), .ip2(\cache_tag[12][21] ), .op(n12183) );
  nand2_1 U14928 ( .ip1(n12179), .ip2(\cache_tag[6][21] ), .op(n12182) );
  nand2_1 U14929 ( .ip1(n12233), .ip2(\cache_tag[0][21] ), .op(n12181) );
  nand2_1 U14930 ( .ip1(n12235), .ip2(\cache_tag[10][21] ), .op(n12180) );
  nand4_1 U14931 ( .ip1(n12183), .ip2(n12182), .ip3(n12181), .ip4(n12180), 
        .op(n12184) );
  nor4_1 U14932 ( .ip1(n12187), .ip2(n12186), .ip3(n12185), .ip4(n12184), .op(
        n12188) );
  nor2_1 U14933 ( .ip1(n12188), .ip2(n12252), .op(n12190) );
  and2_1 U14934 ( .ip1(n12254), .ip2(addr_resp[29]), .op(n12189) );
  ab_or_c_or_d U14935 ( .ip1(addr_mem[29]), .ip2(n12257), .ip3(n12190), .ip4(
        n12189), .op(n4754) );
  nand2_1 U14936 ( .ip1(n9669), .ip2(\cache_tag[11][22] ), .op(n12195) );
  nand2_1 U14937 ( .ip1(n12240), .ip2(\cache_tag[5][22] ), .op(n12194) );
  nand2_1 U14938 ( .ip1(n12242), .ip2(\cache_tag[13][22] ), .op(n12193) );
  nand2_1 U14939 ( .ip1(n12191), .ip2(\cache_tag[8][22] ), .op(n12192) );
  nand4_1 U14940 ( .ip1(n12195), .ip2(n12194), .ip3(n12193), .ip4(n12192), 
        .op(n12215) );
  nand2_1 U14941 ( .ip1(n12220), .ip2(\cache_tag[14][22] ), .op(n12200) );
  nand2_1 U14942 ( .ip1(n12233), .ip2(\cache_tag[0][22] ), .op(n12199) );
  nand2_1 U14943 ( .ip1(n12196), .ip2(\cache_tag[10][22] ), .op(n12198) );
  nand2_1 U14944 ( .ip1(n12241), .ip2(\cache_tag[9][22] ), .op(n12197) );
  nand4_1 U14945 ( .ip1(n12200), .ip2(n12199), .ip3(n12198), .ip4(n12197), 
        .op(n12214) );
  nand2_1 U14946 ( .ip1(n12201), .ip2(\cache_tag[4][22] ), .op(n12206) );
  nand2_1 U14947 ( .ip1(n12219), .ip2(\cache_tag[3][22] ), .op(n12205) );
  nand2_1 U14948 ( .ip1(n12228), .ip2(\cache_tag[2][22] ), .op(n12204) );
  nand2_1 U14949 ( .ip1(n12202), .ip2(\cache_tag[7][22] ), .op(n12203) );
  nand4_1 U14950 ( .ip1(n12206), .ip2(n12205), .ip3(n12204), .ip4(n12203), 
        .op(n12213) );
  nand2_1 U14951 ( .ip1(n12207), .ip2(\cache_tag[12][22] ), .op(n12211) );
  nand2_1 U14952 ( .ip1(n10305), .ip2(\cache_tag[6][22] ), .op(n12210) );
  nand2_1 U14953 ( .ip1(n11979), .ip2(\cache_tag[1][22] ), .op(n12209) );
  nand2_1 U14954 ( .ip1(n12221), .ip2(\cache_tag[15][22] ), .op(n12208) );
  nand4_1 U14955 ( .ip1(n12211), .ip2(n12210), .ip3(n12209), .ip4(n12208), 
        .op(n12212) );
  nor4_1 U14956 ( .ip1(n12215), .ip2(n12214), .ip3(n12213), .ip4(n12212), .op(
        n12216) );
  nor2_1 U14957 ( .ip1(n12216), .ip2(n12252), .op(n12218) );
  and2_1 U14958 ( .ip1(n12254), .ip2(addr_resp[30]), .op(n12217) );
  ab_or_c_or_d U14959 ( .ip1(addr_mem[30]), .ip2(n12257), .ip3(n12218), .ip4(
        n12217), .op(n4753) );
  nand2_1 U14960 ( .ip1(n12219), .ip2(\cache_tag[3][23] ), .op(n12225) );
  nand2_1 U14961 ( .ip1(n12220), .ip2(\cache_tag[14][23] ), .op(n12224) );
  nand2_1 U14962 ( .ip1(n12221), .ip2(\cache_tag[15][23] ), .op(n12223) );
  nand2_1 U14963 ( .ip1(n11943), .ip2(\cache_tag[1][23] ), .op(n12222) );
  nand4_1 U14964 ( .ip1(n12225), .ip2(n12224), .ip3(n12223), .ip4(n12222), 
        .op(n12251) );
  nand2_1 U14965 ( .ip1(n12226), .ip2(\cache_tag[7][23] ), .op(n12232) );
  nand2_1 U14966 ( .ip1(n12227), .ip2(\cache_tag[12][23] ), .op(n12231) );
  nand2_1 U14967 ( .ip1(n12228), .ip2(\cache_tag[2][23] ), .op(n12230) );
  nand2_1 U14968 ( .ip1(n9669), .ip2(\cache_tag[11][23] ), .op(n12229) );
  nand4_1 U14969 ( .ip1(n12232), .ip2(n12231), .ip3(n12230), .ip4(n12229), 
        .op(n12250) );
  nand2_1 U14970 ( .ip1(n12233), .ip2(\cache_tag[0][23] ), .op(n12239) );
  nand2_1 U14971 ( .ip1(n10305), .ip2(\cache_tag[6][23] ), .op(n12238) );
  nand2_1 U14972 ( .ip1(n12234), .ip2(\cache_tag[8][23] ), .op(n12237) );
  nand2_1 U14973 ( .ip1(n12235), .ip2(\cache_tag[10][23] ), .op(n12236) );
  nand4_1 U14974 ( .ip1(n12239), .ip2(n12238), .ip3(n12237), .ip4(n12236), 
        .op(n12249) );
  nand2_1 U14975 ( .ip1(n12240), .ip2(\cache_tag[5][23] ), .op(n12247) );
  nand2_1 U14976 ( .ip1(n12241), .ip2(\cache_tag[9][23] ), .op(n12246) );
  nand2_1 U14977 ( .ip1(n12242), .ip2(\cache_tag[13][23] ), .op(n12245) );
  nand2_1 U14978 ( .ip1(n12243), .ip2(\cache_tag[4][23] ), .op(n12244) );
  nand4_1 U14979 ( .ip1(n12247), .ip2(n12246), .ip3(n12245), .ip4(n12244), 
        .op(n12248) );
  nor4_1 U14980 ( .ip1(n12251), .ip2(n12250), .ip3(n12249), .ip4(n12248), .op(
        n12253) );
  nor2_1 U14981 ( .ip1(n12253), .ip2(n12252), .op(n12256) );
  and2_1 U14982 ( .ip1(n12254), .ip2(addr_resp[31]), .op(n12255) );
  ab_or_c_or_d U14983 ( .ip1(addr_mem[31]), .ip2(n12257), .ip3(n12256), .ip4(
        n12255), .op(n4752) );
  nand2_1 U14985 ( .ip1(n12261), .ip2(cache_miss_count[29]), .op(n12259) );
  inv_1 U14986 ( .ip(cache_miss_count[30]), .op(n12260) );
  nor2_1 U14987 ( .ip1(n12259), .ip2(n12260), .op(n12258) );
  xor2_1 U14988 ( .ip1(n12258), .ip2(cache_miss_count[31]), .op(n4750) );
  mux2_1 U14989 ( .ip1(n12260), .ip2(cache_miss_count[30]), .s(n12259), .op(
        n4749) );
  xor2_1 U14990 ( .ip1(n12261), .ip2(cache_miss_count[29]), .op(n4748) );
  xor2_1 U14991 ( .ip1(n12262), .ip2(cache_miss_count[27]), .op(n4746) );
  xor2_1 U14992 ( .ip1(n12263), .ip2(cache_miss_count[25]), .op(n4744) );
  xor2_1 U14993 ( .ip1(n12264), .ip2(cache_miss_count[23]), .op(n4742) );
  xor2_1 U14994 ( .ip1(n12265), .ip2(cache_miss_count[21]), .op(n4740) );
  xor2_1 U14995 ( .ip1(n12266), .ip2(cache_miss_count[19]), .op(n4738) );
  inv_1 U14996 ( .ip(cache_miss_count[18]), .op(n12268) );
  and2_1 U14997 ( .ip1(cache_miss_count[16]), .ip2(n12270), .op(n12272) );
  nand2_1 U14998 ( .ip1(cache_miss_count[17]), .ip2(n12272), .op(n12267) );
  mux2_1 U14999 ( .ip1(n12268), .ip2(cache_miss_count[18]), .s(n12267), .op(
        n4737) );
  inv_1 U15000 ( .ip(cache_miss_count[17]), .op(n12269) );
  mux2_1 U15001 ( .ip1(cache_miss_count[17]), .ip2(n12269), .s(n12272), .op(
        n4736) );
  nor2_1 U15002 ( .ip1(cache_miss_count[16]), .ip2(n12270), .op(n12271) );
  nor2_1 U15003 ( .ip1(n12272), .ip2(n12271), .op(n4735) );
  inv_1 U15004 ( .ip(cache_miss_count[14]), .op(n12274) );
  mux2_1 U15005 ( .ip1(cache_miss_count[14]), .ip2(n12274), .s(n12273), .op(
        n4733) );
  inv_1 U15006 ( .ip(cache_miss_count[12]), .op(n12276) );
  mux2_1 U15007 ( .ip1(cache_miss_count[12]), .ip2(n12276), .s(n12275), .op(
        n4731) );
  inv_1 U15008 ( .ip(cache_miss_count[10]), .op(n12278) );
  mux2_1 U15009 ( .ip1(cache_miss_count[10]), .ip2(n12278), .s(n12277), .op(
        n4729) );
  inv_1 U15010 ( .ip(cache_miss_count[8]), .op(n12280) );
  mux2_1 U15011 ( .ip1(cache_miss_count[8]), .ip2(n12280), .s(n12279), .op(
        n4727) );
  inv_1 U15012 ( .ip(n12281), .op(n12284) );
  nor2_1 U15013 ( .ip1(n12282), .ip2(cache_miss_count[6]), .op(n12283) );
  nor2_1 U15014 ( .ip1(n12284), .ip2(n12283), .op(n4725) );
  xor2_1 U15015 ( .ip1(n12285), .ip2(cache_miss_count[4]), .op(n4723) );
  xor2_1 U15016 ( .ip1(n12286), .ip2(cache_miss_count[2]), .op(n4721) );
  inv_1 U15017 ( .ip(cache_miss_count[0]), .op(n12289) );
  nand2_1 U15018 ( .ip1(n12287), .ip2(miss), .op(n12288) );
  mux2_1 U15019 ( .ip1(n12289), .ip2(cache_miss_count[0]), .s(n12288), .op(
        n4719) );
  nand2_1 U15020 ( .ip1(n12293), .ip2(cache_hit_count[29]), .op(n12291) );
  inv_1 U15021 ( .ip(cache_hit_count[30]), .op(n12292) );
  nor2_1 U15022 ( .ip1(n12291), .ip2(n12292), .op(n12290) );
  xor2_1 U15023 ( .ip1(n12290), .ip2(cache_hit_count[31]), .op(n4718) );
  mux2_1 U15024 ( .ip1(n12292), .ip2(cache_hit_count[30]), .s(n12291), .op(
        n4717) );
  xor2_1 U15025 ( .ip1(n12293), .ip2(cache_hit_count[29]), .op(n4716) );
  xor2_1 U15026 ( .ip1(n12294), .ip2(cache_hit_count[27]), .op(n4714) );
  xor2_1 U15027 ( .ip1(n12295), .ip2(cache_hit_count[25]), .op(n4712) );
  xor2_1 U15028 ( .ip1(n12296), .ip2(cache_hit_count[23]), .op(n4710) );
  inv_1 U15029 ( .ip(n12297), .op(n12301) );
  nor2_1 U15030 ( .ip1(n12299), .ip2(n12298), .op(n12304) );
  nor2_1 U15031 ( .ip1(cache_hit_count[21]), .ip2(n12304), .op(n12300) );
  nor2_1 U15032 ( .ip1(n12301), .ip2(n12300), .op(n4708) );
  nor2_1 U15033 ( .ip1(cache_hit_count[20]), .ip2(n12302), .op(n12303) );
  nor2_1 U15034 ( .ip1(n12304), .ip2(n12303), .op(n4707) );
  inv_1 U15035 ( .ip(cache_hit_count[18]), .op(n12306) );
  mux2_1 U15036 ( .ip1(cache_hit_count[18]), .ip2(n12306), .s(n12305), .op(
        n4705) );
  inv_1 U15037 ( .ip(n12307), .op(n12310) );
  nor2_1 U15038 ( .ip1(n12308), .ip2(cache_hit_count[16]), .op(n12309) );
  nor2_1 U15039 ( .ip1(n12310), .ip2(n12309), .op(n4703) );
  xor2_1 U15040 ( .ip1(n12311), .ip2(cache_hit_count[14]), .op(n4701) );
  mux2_1 U15041 ( .ip1(cache_hit_count[11]), .ip2(n12313), .s(n12312), .op(
        n4698) );
  mux2_1 U15042 ( .ip1(cache_hit_count[9]), .ip2(n12315), .s(n12314), .op(
        n4696) );
  inv_1 U15043 ( .ip(n12317), .op(n12316) );
  mux2_1 U15044 ( .ip1(n12317), .ip2(n12316), .s(cache_hit_count[7]), .op(
        n4694) );
  xor2_1 U15045 ( .ip1(n12318), .ip2(cache_hit_count[5]), .op(n4692) );
  xor2_1 U15046 ( .ip1(n12319), .ip2(cache_hit_count[3]), .op(n4690) );
  xor2_1 U15047 ( .ip1(n12320), .ip2(cache_hit_count[1]), .op(n4688) );
  inv_1 U15048 ( .ip(N3615), .op(n127) );
  inv_1 U15049 ( .ip(N3612), .op(n125) );
  inv_1 U15050 ( .ip(N3609), .op(n123) );
  inv_1 U15051 ( .ip(N3606), .op(n121) );
  inv_1 U15052 ( .ip(N3603), .op(n119) );
  inv_1 U15053 ( .ip(N3600), .op(n117) );
  inv_1 U15054 ( .ip(N3597), .op(n115) );
  inv_1 U15055 ( .ip(N3594), .op(n113) );
  inv_1 U15056 ( .ip(N3591), .op(n111) );
  inv_1 U15057 ( .ip(N3588), .op(n109) );
  inv_1 U15058 ( .ip(N3585), .op(n107) );
  inv_1 U15059 ( .ip(N3582), .op(n105) );
  inv_1 U15060 ( .ip(N3579), .op(n103) );
  inv_1 U15061 ( .ip(N3576), .op(n101) );
  inv_1 U15062 ( .ip(N3573), .op(n99) );
  inv_1 U15063 ( .ip(N3570), .op(n97) );
  inv_1 U15064 ( .ip(N3567), .op(n95) );
  inv_1 U15065 ( .ip(N3564), .op(n93) );
  inv_1 U15066 ( .ip(N3561), .op(n91) );
  inv_1 U15067 ( .ip(N3558), .op(n89) );
  inv_1 U15068 ( .ip(N3555), .op(n87) );
  inv_1 U15069 ( .ip(N3552), .op(n85) );
  inv_1 U15070 ( .ip(N3549), .op(n83) );
  inv_1 U15071 ( .ip(N3546), .op(n81) );
  inv_1 U15072 ( .ip(N3543), .op(n79) );
  inv_1 U15073 ( .ip(N3540), .op(n77) );
  inv_1 U15074 ( .ip(N3537), .op(n75) );
  inv_1 U15075 ( .ip(N3534), .op(n73) );
  inv_1 U15076 ( .ip(N3531), .op(n71) );
  inv_1 U15077 ( .ip(N3528), .op(n69) );
  inv_1 U15078 ( .ip(N3525), .op(n67) );
  inv_1 U15079 ( .ip(N3522), .op(n65) );
  inv_1 U15080 ( .ip(N3519), .op(n63) );
  inv_1 U15081 ( .ip(N3516), .op(n61) );
  inv_1 U15082 ( .ip(N3513), .op(n59) );
  inv_1 U15083 ( .ip(N3510), .op(n57) );
  inv_1 U15084 ( .ip(N3507), .op(n55) );
  inv_1 U15085 ( .ip(N3504), .op(n53) );
  inv_1 U15086 ( .ip(N3501), .op(n51) );
  inv_1 U15087 ( .ip(N3498), .op(n49) );
  inv_1 U15088 ( .ip(N3495), .op(n47) );
  inv_1 U15089 ( .ip(N3492), .op(n45) );
  inv_1 U15090 ( .ip(N3489), .op(n43) );
  inv_1 U15091 ( .ip(N3486), .op(n41) );
  inv_1 U15092 ( .ip(N3483), .op(n39) );
  inv_1 U15093 ( .ip(N3480), .op(n37) );
  inv_1 U15094 ( .ip(N3477), .op(n35) );
  inv_1 U15095 ( .ip(N3474), .op(n33) );
  inv_1 U15096 ( .ip(N3471), .op(n31) );
  inv_1 U15097 ( .ip(N3468), .op(n29) );
  inv_1 U15098 ( .ip(N3465), .op(n27) );
  inv_1 U15099 ( .ip(N3462), .op(n25) );
  inv_1 U15100 ( .ip(N3459), .op(n23) );
  inv_1 U15101 ( .ip(N3456), .op(n21) );
  inv_1 U15102 ( .ip(N3453), .op(n19) );
  inv_1 U15103 ( .ip(N3450), .op(n17) );
  inv_1 U15104 ( .ip(N3447), .op(n15) );
  inv_1 U15105 ( .ip(N3444), .op(n13) );
  inv_1 U15106 ( .ip(N3441), .op(n11) );
  inv_1 U15107 ( .ip(N3438), .op(n9) );
  inv_1 U15108 ( .ip(N3435), .op(n7) );
  inv_1 U15109 ( .ip(N3432), .op(n5) );
  inv_1 U15110 ( .ip(N3429), .op(n3) );
  inv_1 U15111 ( .ip(N3426), .op(n1) );
endmodule

