
module CacheController ( rst, clk, wr, rd, data_rd, data_wr, addr_req, 
        addr_resp, rdy, busy, wr_mem, rd_mem, busy_mem, data_rd_mem, 
        data_wr_mem, addr_mem, cache_miss_count, cache_hit_count );
  output [31:0] data_rd;
  input [31:0] data_wr;
  input [31:0] addr_req;
  output [31:0] addr_resp;
  input [31:0] data_rd_mem;
  output [31:0] data_wr_mem;
  output [31:0] addr_mem;
  output [31:0] cache_miss_count;
  output [31:0] cache_hit_count;
  input rst, clk, wr, rd, busy_mem;
  output rdy, busy, wr_mem, rd_mem;
  wire   valid, dirty, miss, mem_done, hit, \cache_tag_A[7][24] ,
         \cache_tag_A[7][23] , \cache_tag_A[7][22] , \cache_tag_A[7][21] ,
         \cache_tag_A[7][20] , \cache_tag_A[7][19] , \cache_tag_A[7][18] ,
         \cache_tag_A[7][17] , \cache_tag_A[7][16] , \cache_tag_A[7][15] ,
         \cache_tag_A[7][14] , \cache_tag_A[7][13] , \cache_tag_A[7][12] ,
         \cache_tag_A[7][11] , \cache_tag_A[7][10] , \cache_tag_A[7][9] ,
         \cache_tag_A[7][8] , \cache_tag_A[7][7] , \cache_tag_A[7][6] ,
         \cache_tag_A[7][5] , \cache_tag_A[7][4] , \cache_tag_A[7][3] ,
         \cache_tag_A[7][2] , \cache_tag_A[7][1] , \cache_tag_A[7][0] ,
         \cache_tag_A[6][24] , \cache_tag_A[6][23] , \cache_tag_A[6][22] ,
         \cache_tag_A[6][21] , \cache_tag_A[6][20] , \cache_tag_A[6][19] ,
         \cache_tag_A[6][18] , \cache_tag_A[6][17] , \cache_tag_A[6][16] ,
         \cache_tag_A[6][15] , \cache_tag_A[6][14] , \cache_tag_A[6][13] ,
         \cache_tag_A[6][12] , \cache_tag_A[6][11] , \cache_tag_A[6][10] ,
         \cache_tag_A[6][9] , \cache_tag_A[6][8] , \cache_tag_A[6][7] ,
         \cache_tag_A[6][6] , \cache_tag_A[6][5] , \cache_tag_A[6][4] ,
         \cache_tag_A[6][3] , \cache_tag_A[6][2] , \cache_tag_A[6][1] ,
         \cache_tag_A[6][0] , \cache_tag_A[5][24] , \cache_tag_A[5][23] ,
         \cache_tag_A[5][22] , \cache_tag_A[5][21] , \cache_tag_A[5][20] ,
         \cache_tag_A[5][19] , \cache_tag_A[5][18] , \cache_tag_A[5][17] ,
         \cache_tag_A[5][16] , \cache_tag_A[5][15] , \cache_tag_A[5][14] ,
         \cache_tag_A[5][13] , \cache_tag_A[5][12] , \cache_tag_A[5][11] ,
         \cache_tag_A[5][10] , \cache_tag_A[5][9] , \cache_tag_A[5][8] ,
         \cache_tag_A[5][7] , \cache_tag_A[5][6] , \cache_tag_A[5][5] ,
         \cache_tag_A[5][4] , \cache_tag_A[5][3] , \cache_tag_A[5][2] ,
         \cache_tag_A[5][1] , \cache_tag_A[5][0] , \cache_tag_A[4][24] ,
         \cache_tag_A[4][23] , \cache_tag_A[4][22] , \cache_tag_A[4][21] ,
         \cache_tag_A[4][20] , \cache_tag_A[4][19] , \cache_tag_A[4][18] ,
         \cache_tag_A[4][17] , \cache_tag_A[4][16] , \cache_tag_A[4][15] ,
         \cache_tag_A[4][14] , \cache_tag_A[4][13] , \cache_tag_A[4][12] ,
         \cache_tag_A[4][11] , \cache_tag_A[4][10] , \cache_tag_A[4][9] ,
         \cache_tag_A[4][8] , \cache_tag_A[4][7] , \cache_tag_A[4][6] ,
         \cache_tag_A[4][5] , \cache_tag_A[4][4] , \cache_tag_A[4][3] ,
         \cache_tag_A[4][2] , \cache_tag_A[4][1] , \cache_tag_A[4][0] ,
         \cache_tag_A[3][24] , \cache_tag_A[3][23] , \cache_tag_A[3][22] ,
         \cache_tag_A[3][21] , \cache_tag_A[3][20] , \cache_tag_A[3][19] ,
         \cache_tag_A[3][18] , \cache_tag_A[3][17] , \cache_tag_A[3][16] ,
         \cache_tag_A[3][15] , \cache_tag_A[3][14] , \cache_tag_A[3][13] ,
         \cache_tag_A[3][12] , \cache_tag_A[3][11] , \cache_tag_A[3][10] ,
         \cache_tag_A[3][9] , \cache_tag_A[3][8] , \cache_tag_A[3][7] ,
         \cache_tag_A[3][6] , \cache_tag_A[3][5] , \cache_tag_A[3][4] ,
         \cache_tag_A[3][3] , \cache_tag_A[3][2] , \cache_tag_A[3][1] ,
         \cache_tag_A[3][0] , \cache_tag_A[2][24] , \cache_tag_A[2][23] ,
         \cache_tag_A[2][22] , \cache_tag_A[2][21] , \cache_tag_A[2][20] ,
         \cache_tag_A[2][19] , \cache_tag_A[2][18] , \cache_tag_A[2][17] ,
         \cache_tag_A[2][16] , \cache_tag_A[2][15] , \cache_tag_A[2][14] ,
         \cache_tag_A[2][13] , \cache_tag_A[2][12] , \cache_tag_A[2][11] ,
         \cache_tag_A[2][10] , \cache_tag_A[2][9] , \cache_tag_A[2][8] ,
         \cache_tag_A[2][7] , \cache_tag_A[2][6] , \cache_tag_A[2][5] ,
         \cache_tag_A[2][4] , \cache_tag_A[2][3] , \cache_tag_A[2][2] ,
         \cache_tag_A[2][1] , \cache_tag_A[2][0] , \cache_tag_A[1][24] ,
         \cache_tag_A[1][23] , \cache_tag_A[1][22] , \cache_tag_A[1][21] ,
         \cache_tag_A[1][20] , \cache_tag_A[1][19] , \cache_tag_A[1][18] ,
         \cache_tag_A[1][17] , \cache_tag_A[1][16] , \cache_tag_A[1][15] ,
         \cache_tag_A[1][14] , \cache_tag_A[1][13] , \cache_tag_A[1][12] ,
         \cache_tag_A[1][11] , \cache_tag_A[1][10] , \cache_tag_A[1][9] ,
         \cache_tag_A[1][8] , \cache_tag_A[1][7] , \cache_tag_A[1][6] ,
         \cache_tag_A[1][5] , \cache_tag_A[1][4] , \cache_tag_A[1][3] ,
         \cache_tag_A[1][2] , \cache_tag_A[1][1] , \cache_tag_A[1][0] ,
         \cache_tag_A[0][24] , \cache_tag_A[0][23] , \cache_tag_A[0][22] ,
         \cache_tag_A[0][21] , \cache_tag_A[0][20] , \cache_tag_A[0][19] ,
         \cache_tag_A[0][18] , \cache_tag_A[0][17] , \cache_tag_A[0][16] ,
         \cache_tag_A[0][15] , \cache_tag_A[0][14] , \cache_tag_A[0][13] ,
         \cache_tag_A[0][12] , \cache_tag_A[0][11] , \cache_tag_A[0][10] ,
         \cache_tag_A[0][9] , \cache_tag_A[0][8] , \cache_tag_A[0][7] ,
         \cache_tag_A[0][6] , \cache_tag_A[0][5] , \cache_tag_A[0][4] ,
         \cache_tag_A[0][3] , \cache_tag_A[0][2] , \cache_tag_A[0][1] ,
         \cache_tag_A[0][0] , \cache_data_A[7][127] , \cache_data_A[7][126] ,
         \cache_data_A[7][125] , \cache_data_A[7][124] ,
         \cache_data_A[7][123] , \cache_data_A[7][122] ,
         \cache_data_A[7][121] , \cache_data_A[7][120] ,
         \cache_data_A[7][119] , \cache_data_A[7][118] ,
         \cache_data_A[7][117] , \cache_data_A[7][116] ,
         \cache_data_A[7][115] , \cache_data_A[7][114] ,
         \cache_data_A[7][113] , \cache_data_A[7][112] ,
         \cache_data_A[7][111] , \cache_data_A[7][110] ,
         \cache_data_A[7][109] , \cache_data_A[7][108] ,
         \cache_data_A[7][107] , \cache_data_A[7][106] ,
         \cache_data_A[7][105] , \cache_data_A[7][104] ,
         \cache_data_A[7][103] , \cache_data_A[7][102] ,
         \cache_data_A[7][101] , \cache_data_A[7][100] , \cache_data_A[7][99] ,
         \cache_data_A[7][98] , \cache_data_A[7][97] , \cache_data_A[7][96] ,
         \cache_data_A[7][95] , \cache_data_A[7][94] , \cache_data_A[7][93] ,
         \cache_data_A[7][92] , \cache_data_A[7][91] , \cache_data_A[7][90] ,
         \cache_data_A[7][89] , \cache_data_A[7][88] , \cache_data_A[7][87] ,
         \cache_data_A[7][86] , \cache_data_A[7][85] , \cache_data_A[7][84] ,
         \cache_data_A[7][83] , \cache_data_A[7][82] , \cache_data_A[7][81] ,
         \cache_data_A[7][80] , \cache_data_A[7][79] , \cache_data_A[7][78] ,
         \cache_data_A[7][77] , \cache_data_A[7][76] , \cache_data_A[7][75] ,
         \cache_data_A[7][74] , \cache_data_A[7][73] , \cache_data_A[7][72] ,
         \cache_data_A[7][71] , \cache_data_A[7][70] , \cache_data_A[7][69] ,
         \cache_data_A[7][68] , \cache_data_A[7][67] , \cache_data_A[7][66] ,
         \cache_data_A[7][65] , \cache_data_A[7][64] , \cache_data_A[7][63] ,
         \cache_data_A[7][62] , \cache_data_A[7][61] , \cache_data_A[7][60] ,
         \cache_data_A[7][59] , \cache_data_A[7][58] , \cache_data_A[7][57] ,
         \cache_data_A[7][56] , \cache_data_A[7][55] , \cache_data_A[7][54] ,
         \cache_data_A[7][53] , \cache_data_A[7][52] , \cache_data_A[7][51] ,
         \cache_data_A[7][50] , \cache_data_A[7][49] , \cache_data_A[7][48] ,
         \cache_data_A[7][47] , \cache_data_A[7][46] , \cache_data_A[7][45] ,
         \cache_data_A[7][44] , \cache_data_A[7][43] , \cache_data_A[7][42] ,
         \cache_data_A[7][41] , \cache_data_A[7][40] , \cache_data_A[7][39] ,
         \cache_data_A[7][38] , \cache_data_A[7][37] , \cache_data_A[7][36] ,
         \cache_data_A[7][35] , \cache_data_A[7][34] , \cache_data_A[7][33] ,
         \cache_data_A[7][32] , \cache_data_A[7][31] , \cache_data_A[7][30] ,
         \cache_data_A[7][29] , \cache_data_A[7][28] , \cache_data_A[7][27] ,
         \cache_data_A[7][26] , \cache_data_A[7][25] , \cache_data_A[7][24] ,
         \cache_data_A[7][23] , \cache_data_A[7][22] , \cache_data_A[7][21] ,
         \cache_data_A[7][20] , \cache_data_A[7][19] , \cache_data_A[7][18] ,
         \cache_data_A[7][17] , \cache_data_A[7][16] , \cache_data_A[7][15] ,
         \cache_data_A[7][14] , \cache_data_A[7][13] , \cache_data_A[7][12] ,
         \cache_data_A[7][11] , \cache_data_A[7][10] , \cache_data_A[7][9] ,
         \cache_data_A[7][8] , \cache_data_A[7][7] , \cache_data_A[7][6] ,
         \cache_data_A[7][5] , \cache_data_A[7][4] , \cache_data_A[7][3] ,
         \cache_data_A[7][2] , \cache_data_A[7][1] , \cache_data_A[7][0] ,
         \cache_data_A[6][127] , \cache_data_A[6][126] ,
         \cache_data_A[6][125] , \cache_data_A[6][124] ,
         \cache_data_A[6][123] , \cache_data_A[6][122] ,
         \cache_data_A[6][121] , \cache_data_A[6][120] ,
         \cache_data_A[6][119] , \cache_data_A[6][118] ,
         \cache_data_A[6][117] , \cache_data_A[6][116] ,
         \cache_data_A[6][115] , \cache_data_A[6][114] ,
         \cache_data_A[6][113] , \cache_data_A[6][112] ,
         \cache_data_A[6][111] , \cache_data_A[6][110] ,
         \cache_data_A[6][109] , \cache_data_A[6][108] ,
         \cache_data_A[6][107] , \cache_data_A[6][106] ,
         \cache_data_A[6][105] , \cache_data_A[6][104] ,
         \cache_data_A[6][103] , \cache_data_A[6][102] ,
         \cache_data_A[6][101] , \cache_data_A[6][100] , \cache_data_A[6][99] ,
         \cache_data_A[6][98] , \cache_data_A[6][97] , \cache_data_A[6][96] ,
         \cache_data_A[6][95] , \cache_data_A[6][94] , \cache_data_A[6][93] ,
         \cache_data_A[6][92] , \cache_data_A[6][91] , \cache_data_A[6][90] ,
         \cache_data_A[6][89] , \cache_data_A[6][88] , \cache_data_A[6][87] ,
         \cache_data_A[6][86] , \cache_data_A[6][85] , \cache_data_A[6][84] ,
         \cache_data_A[6][83] , \cache_data_A[6][82] , \cache_data_A[6][81] ,
         \cache_data_A[6][80] , \cache_data_A[6][79] , \cache_data_A[6][78] ,
         \cache_data_A[6][77] , \cache_data_A[6][76] , \cache_data_A[6][75] ,
         \cache_data_A[6][74] , \cache_data_A[6][73] , \cache_data_A[6][72] ,
         \cache_data_A[6][71] , \cache_data_A[6][70] , \cache_data_A[6][69] ,
         \cache_data_A[6][68] , \cache_data_A[6][67] , \cache_data_A[6][66] ,
         \cache_data_A[6][65] , \cache_data_A[6][64] , \cache_data_A[6][63] ,
         \cache_data_A[6][62] , \cache_data_A[6][61] , \cache_data_A[6][60] ,
         \cache_data_A[6][59] , \cache_data_A[6][58] , \cache_data_A[6][57] ,
         \cache_data_A[6][56] , \cache_data_A[6][55] , \cache_data_A[6][54] ,
         \cache_data_A[6][53] , \cache_data_A[6][52] , \cache_data_A[6][51] ,
         \cache_data_A[6][50] , \cache_data_A[6][49] , \cache_data_A[6][48] ,
         \cache_data_A[6][47] , \cache_data_A[6][46] , \cache_data_A[6][45] ,
         \cache_data_A[6][44] , \cache_data_A[6][43] , \cache_data_A[6][42] ,
         \cache_data_A[6][41] , \cache_data_A[6][40] , \cache_data_A[6][39] ,
         \cache_data_A[6][38] , \cache_data_A[6][37] , \cache_data_A[6][36] ,
         \cache_data_A[6][35] , \cache_data_A[6][34] , \cache_data_A[6][33] ,
         \cache_data_A[6][32] , \cache_data_A[6][31] , \cache_data_A[6][30] ,
         \cache_data_A[6][29] , \cache_data_A[6][28] , \cache_data_A[6][27] ,
         \cache_data_A[6][26] , \cache_data_A[6][25] , \cache_data_A[6][24] ,
         \cache_data_A[6][23] , \cache_data_A[6][22] , \cache_data_A[6][21] ,
         \cache_data_A[6][20] , \cache_data_A[6][19] , \cache_data_A[6][18] ,
         \cache_data_A[6][17] , \cache_data_A[6][16] , \cache_data_A[6][15] ,
         \cache_data_A[6][14] , \cache_data_A[6][13] , \cache_data_A[6][12] ,
         \cache_data_A[6][11] , \cache_data_A[6][10] , \cache_data_A[6][9] ,
         \cache_data_A[6][8] , \cache_data_A[6][7] , \cache_data_A[6][6] ,
         \cache_data_A[6][5] , \cache_data_A[6][4] , \cache_data_A[6][3] ,
         \cache_data_A[6][2] , \cache_data_A[6][1] , \cache_data_A[6][0] ,
         \cache_data_A[5][127] , \cache_data_A[5][126] ,
         \cache_data_A[5][125] , \cache_data_A[5][124] ,
         \cache_data_A[5][123] , \cache_data_A[5][122] ,
         \cache_data_A[5][121] , \cache_data_A[5][120] ,
         \cache_data_A[5][119] , \cache_data_A[5][118] ,
         \cache_data_A[5][117] , \cache_data_A[5][116] ,
         \cache_data_A[5][115] , \cache_data_A[5][114] ,
         \cache_data_A[5][113] , \cache_data_A[5][112] ,
         \cache_data_A[5][111] , \cache_data_A[5][110] ,
         \cache_data_A[5][109] , \cache_data_A[5][108] ,
         \cache_data_A[5][107] , \cache_data_A[5][106] ,
         \cache_data_A[5][105] , \cache_data_A[5][104] ,
         \cache_data_A[5][103] , \cache_data_A[5][102] ,
         \cache_data_A[5][101] , \cache_data_A[5][100] , \cache_data_A[5][99] ,
         \cache_data_A[5][98] , \cache_data_A[5][97] , \cache_data_A[5][96] ,
         \cache_data_A[5][95] , \cache_data_A[5][94] , \cache_data_A[5][93] ,
         \cache_data_A[5][92] , \cache_data_A[5][91] , \cache_data_A[5][90] ,
         \cache_data_A[5][89] , \cache_data_A[5][88] , \cache_data_A[5][87] ,
         \cache_data_A[5][86] , \cache_data_A[5][85] , \cache_data_A[5][84] ,
         \cache_data_A[5][83] , \cache_data_A[5][82] , \cache_data_A[5][81] ,
         \cache_data_A[5][80] , \cache_data_A[5][79] , \cache_data_A[5][78] ,
         \cache_data_A[5][77] , \cache_data_A[5][76] , \cache_data_A[5][75] ,
         \cache_data_A[5][74] , \cache_data_A[5][73] , \cache_data_A[5][72] ,
         \cache_data_A[5][71] , \cache_data_A[5][70] , \cache_data_A[5][69] ,
         \cache_data_A[5][68] , \cache_data_A[5][67] , \cache_data_A[5][66] ,
         \cache_data_A[5][65] , \cache_data_A[5][64] , \cache_data_A[5][63] ,
         \cache_data_A[5][62] , \cache_data_A[5][61] , \cache_data_A[5][60] ,
         \cache_data_A[5][59] , \cache_data_A[5][58] , \cache_data_A[5][57] ,
         \cache_data_A[5][56] , \cache_data_A[5][55] , \cache_data_A[5][54] ,
         \cache_data_A[5][53] , \cache_data_A[5][52] , \cache_data_A[5][51] ,
         \cache_data_A[5][50] , \cache_data_A[5][49] , \cache_data_A[5][48] ,
         \cache_data_A[5][47] , \cache_data_A[5][46] , \cache_data_A[5][45] ,
         \cache_data_A[5][44] , \cache_data_A[5][43] , \cache_data_A[5][42] ,
         \cache_data_A[5][41] , \cache_data_A[5][40] , \cache_data_A[5][39] ,
         \cache_data_A[5][38] , \cache_data_A[5][37] , \cache_data_A[5][36] ,
         \cache_data_A[5][35] , \cache_data_A[5][34] , \cache_data_A[5][33] ,
         \cache_data_A[5][32] , \cache_data_A[5][31] , \cache_data_A[5][30] ,
         \cache_data_A[5][29] , \cache_data_A[5][28] , \cache_data_A[5][27] ,
         \cache_data_A[5][26] , \cache_data_A[5][25] , \cache_data_A[5][24] ,
         \cache_data_A[5][23] , \cache_data_A[5][22] , \cache_data_A[5][21] ,
         \cache_data_A[5][20] , \cache_data_A[5][19] , \cache_data_A[5][18] ,
         \cache_data_A[5][17] , \cache_data_A[5][16] , \cache_data_A[5][15] ,
         \cache_data_A[5][14] , \cache_data_A[5][13] , \cache_data_A[5][12] ,
         \cache_data_A[5][11] , \cache_data_A[5][10] , \cache_data_A[5][9] ,
         \cache_data_A[5][8] , \cache_data_A[5][7] , \cache_data_A[5][6] ,
         \cache_data_A[5][5] , \cache_data_A[5][4] , \cache_data_A[5][3] ,
         \cache_data_A[5][2] , \cache_data_A[5][1] , \cache_data_A[5][0] ,
         \cache_data_A[4][127] , \cache_data_A[4][126] ,
         \cache_data_A[4][125] , \cache_data_A[4][124] ,
         \cache_data_A[4][123] , \cache_data_A[4][122] ,
         \cache_data_A[4][121] , \cache_data_A[4][120] ,
         \cache_data_A[4][119] , \cache_data_A[4][118] ,
         \cache_data_A[4][117] , \cache_data_A[4][116] ,
         \cache_data_A[4][115] , \cache_data_A[4][114] ,
         \cache_data_A[4][113] , \cache_data_A[4][112] ,
         \cache_data_A[4][111] , \cache_data_A[4][110] ,
         \cache_data_A[4][109] , \cache_data_A[4][108] ,
         \cache_data_A[4][107] , \cache_data_A[4][106] ,
         \cache_data_A[4][105] , \cache_data_A[4][104] ,
         \cache_data_A[4][103] , \cache_data_A[4][102] ,
         \cache_data_A[4][101] , \cache_data_A[4][100] , \cache_data_A[4][99] ,
         \cache_data_A[4][98] , \cache_data_A[4][97] , \cache_data_A[4][96] ,
         \cache_data_A[4][95] , \cache_data_A[4][94] , \cache_data_A[4][93] ,
         \cache_data_A[4][92] , \cache_data_A[4][91] , \cache_data_A[4][90] ,
         \cache_data_A[4][89] , \cache_data_A[4][88] , \cache_data_A[4][87] ,
         \cache_data_A[4][86] , \cache_data_A[4][85] , \cache_data_A[4][84] ,
         \cache_data_A[4][83] , \cache_data_A[4][82] , \cache_data_A[4][81] ,
         \cache_data_A[4][80] , \cache_data_A[4][79] , \cache_data_A[4][78] ,
         \cache_data_A[4][77] , \cache_data_A[4][76] , \cache_data_A[4][75] ,
         \cache_data_A[4][74] , \cache_data_A[4][73] , \cache_data_A[4][72] ,
         \cache_data_A[4][71] , \cache_data_A[4][70] , \cache_data_A[4][69] ,
         \cache_data_A[4][68] , \cache_data_A[4][67] , \cache_data_A[4][66] ,
         \cache_data_A[4][65] , \cache_data_A[4][64] , \cache_data_A[4][63] ,
         \cache_data_A[4][62] , \cache_data_A[4][61] , \cache_data_A[4][60] ,
         \cache_data_A[4][59] , \cache_data_A[4][58] , \cache_data_A[4][57] ,
         \cache_data_A[4][56] , \cache_data_A[4][55] , \cache_data_A[4][54] ,
         \cache_data_A[4][53] , \cache_data_A[4][52] , \cache_data_A[4][51] ,
         \cache_data_A[4][50] , \cache_data_A[4][49] , \cache_data_A[4][48] ,
         \cache_data_A[4][47] , \cache_data_A[4][46] , \cache_data_A[4][45] ,
         \cache_data_A[4][44] , \cache_data_A[4][43] , \cache_data_A[4][42] ,
         \cache_data_A[4][41] , \cache_data_A[4][40] , \cache_data_A[4][39] ,
         \cache_data_A[4][38] , \cache_data_A[4][37] , \cache_data_A[4][36] ,
         \cache_data_A[4][35] , \cache_data_A[4][34] , \cache_data_A[4][33] ,
         \cache_data_A[4][32] , \cache_data_A[4][31] , \cache_data_A[4][30] ,
         \cache_data_A[4][29] , \cache_data_A[4][28] , \cache_data_A[4][27] ,
         \cache_data_A[4][26] , \cache_data_A[4][25] , \cache_data_A[4][24] ,
         \cache_data_A[4][23] , \cache_data_A[4][22] , \cache_data_A[4][21] ,
         \cache_data_A[4][20] , \cache_data_A[4][19] , \cache_data_A[4][18] ,
         \cache_data_A[4][17] , \cache_data_A[4][16] , \cache_data_A[4][15] ,
         \cache_data_A[4][14] , \cache_data_A[4][13] , \cache_data_A[4][12] ,
         \cache_data_A[4][11] , \cache_data_A[4][10] , \cache_data_A[4][9] ,
         \cache_data_A[4][8] , \cache_data_A[4][7] , \cache_data_A[4][6] ,
         \cache_data_A[4][5] , \cache_data_A[4][4] , \cache_data_A[4][3] ,
         \cache_data_A[4][2] , \cache_data_A[4][1] , \cache_data_A[4][0] ,
         \cache_data_A[3][127] , \cache_data_A[3][126] ,
         \cache_data_A[3][125] , \cache_data_A[3][124] ,
         \cache_data_A[3][123] , \cache_data_A[3][122] ,
         \cache_data_A[3][121] , \cache_data_A[3][120] ,
         \cache_data_A[3][119] , \cache_data_A[3][118] ,
         \cache_data_A[3][117] , \cache_data_A[3][116] ,
         \cache_data_A[3][115] , \cache_data_A[3][114] ,
         \cache_data_A[3][113] , \cache_data_A[3][112] ,
         \cache_data_A[3][111] , \cache_data_A[3][110] ,
         \cache_data_A[3][109] , \cache_data_A[3][108] ,
         \cache_data_A[3][107] , \cache_data_A[3][106] ,
         \cache_data_A[3][105] , \cache_data_A[3][104] ,
         \cache_data_A[3][103] , \cache_data_A[3][102] ,
         \cache_data_A[3][101] , \cache_data_A[3][100] , \cache_data_A[3][99] ,
         \cache_data_A[3][98] , \cache_data_A[3][97] , \cache_data_A[3][96] ,
         \cache_data_A[3][95] , \cache_data_A[3][94] , \cache_data_A[3][93] ,
         \cache_data_A[3][92] , \cache_data_A[3][91] , \cache_data_A[3][90] ,
         \cache_data_A[3][89] , \cache_data_A[3][88] , \cache_data_A[3][87] ,
         \cache_data_A[3][86] , \cache_data_A[3][85] , \cache_data_A[3][84] ,
         \cache_data_A[3][83] , \cache_data_A[3][82] , \cache_data_A[3][81] ,
         \cache_data_A[3][80] , \cache_data_A[3][79] , \cache_data_A[3][78] ,
         \cache_data_A[3][77] , \cache_data_A[3][76] , \cache_data_A[3][75] ,
         \cache_data_A[3][74] , \cache_data_A[3][73] , \cache_data_A[3][72] ,
         \cache_data_A[3][71] , \cache_data_A[3][70] , \cache_data_A[3][69] ,
         \cache_data_A[3][68] , \cache_data_A[3][67] , \cache_data_A[3][66] ,
         \cache_data_A[3][65] , \cache_data_A[3][64] , \cache_data_A[3][63] ,
         \cache_data_A[3][62] , \cache_data_A[3][61] , \cache_data_A[3][60] ,
         \cache_data_A[3][59] , \cache_data_A[3][58] , \cache_data_A[3][57] ,
         \cache_data_A[3][56] , \cache_data_A[3][55] , \cache_data_A[3][54] ,
         \cache_data_A[3][53] , \cache_data_A[3][52] , \cache_data_A[3][51] ,
         \cache_data_A[3][50] , \cache_data_A[3][49] , \cache_data_A[3][48] ,
         \cache_data_A[3][47] , \cache_data_A[3][46] , \cache_data_A[3][45] ,
         \cache_data_A[3][44] , \cache_data_A[3][43] , \cache_data_A[3][42] ,
         \cache_data_A[3][41] , \cache_data_A[3][40] , \cache_data_A[3][39] ,
         \cache_data_A[3][38] , \cache_data_A[3][37] , \cache_data_A[3][36] ,
         \cache_data_A[3][35] , \cache_data_A[3][34] , \cache_data_A[3][33] ,
         \cache_data_A[3][32] , \cache_data_A[3][31] , \cache_data_A[3][30] ,
         \cache_data_A[3][29] , \cache_data_A[3][28] , \cache_data_A[3][27] ,
         \cache_data_A[3][26] , \cache_data_A[3][25] , \cache_data_A[3][24] ,
         \cache_data_A[3][23] , \cache_data_A[3][22] , \cache_data_A[3][21] ,
         \cache_data_A[3][20] , \cache_data_A[3][19] , \cache_data_A[3][18] ,
         \cache_data_A[3][17] , \cache_data_A[3][16] , \cache_data_A[3][15] ,
         \cache_data_A[3][14] , \cache_data_A[3][13] , \cache_data_A[3][12] ,
         \cache_data_A[3][11] , \cache_data_A[3][10] , \cache_data_A[3][9] ,
         \cache_data_A[3][8] , \cache_data_A[3][7] , \cache_data_A[3][6] ,
         \cache_data_A[3][5] , \cache_data_A[3][4] , \cache_data_A[3][3] ,
         \cache_data_A[3][2] , \cache_data_A[3][1] , \cache_data_A[3][0] ,
         \cache_data_A[2][127] , \cache_data_A[2][126] ,
         \cache_data_A[2][125] , \cache_data_A[2][124] ,
         \cache_data_A[2][123] , \cache_data_A[2][122] ,
         \cache_data_A[2][121] , \cache_data_A[2][120] ,
         \cache_data_A[2][119] , \cache_data_A[2][118] ,
         \cache_data_A[2][117] , \cache_data_A[2][116] ,
         \cache_data_A[2][115] , \cache_data_A[2][114] ,
         \cache_data_A[2][113] , \cache_data_A[2][112] ,
         \cache_data_A[2][111] , \cache_data_A[2][110] ,
         \cache_data_A[2][109] , \cache_data_A[2][108] ,
         \cache_data_A[2][107] , \cache_data_A[2][106] ,
         \cache_data_A[2][105] , \cache_data_A[2][104] ,
         \cache_data_A[2][103] , \cache_data_A[2][102] ,
         \cache_data_A[2][101] , \cache_data_A[2][100] , \cache_data_A[2][99] ,
         \cache_data_A[2][98] , \cache_data_A[2][97] , \cache_data_A[2][96] ,
         \cache_data_A[2][95] , \cache_data_A[2][94] , \cache_data_A[2][93] ,
         \cache_data_A[2][92] , \cache_data_A[2][91] , \cache_data_A[2][90] ,
         \cache_data_A[2][89] , \cache_data_A[2][88] , \cache_data_A[2][87] ,
         \cache_data_A[2][86] , \cache_data_A[2][85] , \cache_data_A[2][84] ,
         \cache_data_A[2][83] , \cache_data_A[2][82] , \cache_data_A[2][81] ,
         \cache_data_A[2][80] , \cache_data_A[2][79] , \cache_data_A[2][78] ,
         \cache_data_A[2][77] , \cache_data_A[2][76] , \cache_data_A[2][75] ,
         \cache_data_A[2][74] , \cache_data_A[2][73] , \cache_data_A[2][72] ,
         \cache_data_A[2][71] , \cache_data_A[2][70] , \cache_data_A[2][69] ,
         \cache_data_A[2][68] , \cache_data_A[2][67] , \cache_data_A[2][66] ,
         \cache_data_A[2][65] , \cache_data_A[2][64] , \cache_data_A[2][63] ,
         \cache_data_A[2][62] , \cache_data_A[2][61] , \cache_data_A[2][60] ,
         \cache_data_A[2][59] , \cache_data_A[2][58] , \cache_data_A[2][57] ,
         \cache_data_A[2][56] , \cache_data_A[2][55] , \cache_data_A[2][54] ,
         \cache_data_A[2][53] , \cache_data_A[2][52] , \cache_data_A[2][51] ,
         \cache_data_A[2][50] , \cache_data_A[2][49] , \cache_data_A[2][48] ,
         \cache_data_A[2][47] , \cache_data_A[2][46] , \cache_data_A[2][45] ,
         \cache_data_A[2][44] , \cache_data_A[2][43] , \cache_data_A[2][42] ,
         \cache_data_A[2][41] , \cache_data_A[2][40] , \cache_data_A[2][39] ,
         \cache_data_A[2][38] , \cache_data_A[2][37] , \cache_data_A[2][36] ,
         \cache_data_A[2][35] , \cache_data_A[2][34] , \cache_data_A[2][33] ,
         \cache_data_A[2][32] , \cache_data_A[2][31] , \cache_data_A[2][30] ,
         \cache_data_A[2][29] , \cache_data_A[2][28] , \cache_data_A[2][27] ,
         \cache_data_A[2][26] , \cache_data_A[2][25] , \cache_data_A[2][24] ,
         \cache_data_A[2][23] , \cache_data_A[2][22] , \cache_data_A[2][21] ,
         \cache_data_A[2][20] , \cache_data_A[2][19] , \cache_data_A[2][18] ,
         \cache_data_A[2][17] , \cache_data_A[2][16] , \cache_data_A[2][15] ,
         \cache_data_A[2][14] , \cache_data_A[2][13] , \cache_data_A[2][12] ,
         \cache_data_A[2][11] , \cache_data_A[2][10] , \cache_data_A[2][9] ,
         \cache_data_A[2][8] , \cache_data_A[2][7] , \cache_data_A[2][6] ,
         \cache_data_A[2][5] , \cache_data_A[2][4] , \cache_data_A[2][3] ,
         \cache_data_A[2][2] , \cache_data_A[2][1] , \cache_data_A[2][0] ,
         \cache_data_A[1][127] , \cache_data_A[1][126] ,
         \cache_data_A[1][125] , \cache_data_A[1][124] ,
         \cache_data_A[1][123] , \cache_data_A[1][122] ,
         \cache_data_A[1][121] , \cache_data_A[1][120] ,
         \cache_data_A[1][119] , \cache_data_A[1][118] ,
         \cache_data_A[1][117] , \cache_data_A[1][116] ,
         \cache_data_A[1][115] , \cache_data_A[1][114] ,
         \cache_data_A[1][113] , \cache_data_A[1][112] ,
         \cache_data_A[1][111] , \cache_data_A[1][110] ,
         \cache_data_A[1][109] , \cache_data_A[1][108] ,
         \cache_data_A[1][107] , \cache_data_A[1][106] ,
         \cache_data_A[1][105] , \cache_data_A[1][104] ,
         \cache_data_A[1][103] , \cache_data_A[1][102] ,
         \cache_data_A[1][101] , \cache_data_A[1][100] , \cache_data_A[1][99] ,
         \cache_data_A[1][98] , \cache_data_A[1][97] , \cache_data_A[1][96] ,
         \cache_data_A[1][95] , \cache_data_A[1][94] , \cache_data_A[1][93] ,
         \cache_data_A[1][92] , \cache_data_A[1][91] , \cache_data_A[1][90] ,
         \cache_data_A[1][89] , \cache_data_A[1][88] , \cache_data_A[1][87] ,
         \cache_data_A[1][86] , \cache_data_A[1][85] , \cache_data_A[1][84] ,
         \cache_data_A[1][83] , \cache_data_A[1][82] , \cache_data_A[1][81] ,
         \cache_data_A[1][80] , \cache_data_A[1][79] , \cache_data_A[1][78] ,
         \cache_data_A[1][77] , \cache_data_A[1][76] , \cache_data_A[1][75] ,
         \cache_data_A[1][74] , \cache_data_A[1][73] , \cache_data_A[1][72] ,
         \cache_data_A[1][71] , \cache_data_A[1][70] , \cache_data_A[1][69] ,
         \cache_data_A[1][68] , \cache_data_A[1][67] , \cache_data_A[1][66] ,
         \cache_data_A[1][65] , \cache_data_A[1][64] , \cache_data_A[1][63] ,
         \cache_data_A[1][62] , \cache_data_A[1][61] , \cache_data_A[1][60] ,
         \cache_data_A[1][59] , \cache_data_A[1][58] , \cache_data_A[1][57] ,
         \cache_data_A[1][56] , \cache_data_A[1][55] , \cache_data_A[1][54] ,
         \cache_data_A[1][53] , \cache_data_A[1][52] , \cache_data_A[1][51] ,
         \cache_data_A[1][50] , \cache_data_A[1][49] , \cache_data_A[1][48] ,
         \cache_data_A[1][47] , \cache_data_A[1][46] , \cache_data_A[1][45] ,
         \cache_data_A[1][44] , \cache_data_A[1][43] , \cache_data_A[1][42] ,
         \cache_data_A[1][41] , \cache_data_A[1][40] , \cache_data_A[1][39] ,
         \cache_data_A[1][38] , \cache_data_A[1][37] , \cache_data_A[1][36] ,
         \cache_data_A[1][35] , \cache_data_A[1][34] , \cache_data_A[1][33] ,
         \cache_data_A[1][32] , \cache_data_A[1][31] , \cache_data_A[1][30] ,
         \cache_data_A[1][29] , \cache_data_A[1][28] , \cache_data_A[1][27] ,
         \cache_data_A[1][26] , \cache_data_A[1][25] , \cache_data_A[1][24] ,
         \cache_data_A[1][23] , \cache_data_A[1][22] , \cache_data_A[1][21] ,
         \cache_data_A[1][20] , \cache_data_A[1][19] , \cache_data_A[1][18] ,
         \cache_data_A[1][17] , \cache_data_A[1][16] , \cache_data_A[1][15] ,
         \cache_data_A[1][14] , \cache_data_A[1][13] , \cache_data_A[1][12] ,
         \cache_data_A[1][11] , \cache_data_A[1][10] , \cache_data_A[1][9] ,
         \cache_data_A[1][8] , \cache_data_A[1][7] , \cache_data_A[1][6] ,
         \cache_data_A[1][5] , \cache_data_A[1][4] , \cache_data_A[1][3] ,
         \cache_data_A[1][2] , \cache_data_A[1][1] , \cache_data_A[1][0] ,
         \cache_data_A[0][127] , \cache_data_A[0][126] ,
         \cache_data_A[0][125] , \cache_data_A[0][124] ,
         \cache_data_A[0][123] , \cache_data_A[0][122] ,
         \cache_data_A[0][121] , \cache_data_A[0][120] ,
         \cache_data_A[0][119] , \cache_data_A[0][118] ,
         \cache_data_A[0][117] , \cache_data_A[0][116] ,
         \cache_data_A[0][115] , \cache_data_A[0][114] ,
         \cache_data_A[0][113] , \cache_data_A[0][112] ,
         \cache_data_A[0][111] , \cache_data_A[0][110] ,
         \cache_data_A[0][109] , \cache_data_A[0][108] ,
         \cache_data_A[0][107] , \cache_data_A[0][106] ,
         \cache_data_A[0][105] , \cache_data_A[0][104] ,
         \cache_data_A[0][103] , \cache_data_A[0][102] ,
         \cache_data_A[0][101] , \cache_data_A[0][100] , \cache_data_A[0][99] ,
         \cache_data_A[0][98] , \cache_data_A[0][97] , \cache_data_A[0][96] ,
         \cache_data_A[0][95] , \cache_data_A[0][94] , \cache_data_A[0][93] ,
         \cache_data_A[0][92] , \cache_data_A[0][91] , \cache_data_A[0][90] ,
         \cache_data_A[0][89] , \cache_data_A[0][88] , \cache_data_A[0][87] ,
         \cache_data_A[0][86] , \cache_data_A[0][85] , \cache_data_A[0][84] ,
         \cache_data_A[0][83] , \cache_data_A[0][82] , \cache_data_A[0][81] ,
         \cache_data_A[0][80] , \cache_data_A[0][79] , \cache_data_A[0][78] ,
         \cache_data_A[0][77] , \cache_data_A[0][76] , \cache_data_A[0][75] ,
         \cache_data_A[0][74] , \cache_data_A[0][73] , \cache_data_A[0][72] ,
         \cache_data_A[0][71] , \cache_data_A[0][70] , \cache_data_A[0][69] ,
         \cache_data_A[0][68] , \cache_data_A[0][67] , \cache_data_A[0][66] ,
         \cache_data_A[0][65] , \cache_data_A[0][64] , \cache_data_A[0][63] ,
         \cache_data_A[0][62] , \cache_data_A[0][61] , \cache_data_A[0][60] ,
         \cache_data_A[0][59] , \cache_data_A[0][58] , \cache_data_A[0][57] ,
         \cache_data_A[0][56] , \cache_data_A[0][55] , \cache_data_A[0][54] ,
         \cache_data_A[0][53] , \cache_data_A[0][52] , \cache_data_A[0][51] ,
         \cache_data_A[0][50] , \cache_data_A[0][49] , \cache_data_A[0][48] ,
         \cache_data_A[0][47] , \cache_data_A[0][46] , \cache_data_A[0][45] ,
         \cache_data_A[0][44] , \cache_data_A[0][43] , \cache_data_A[0][42] ,
         \cache_data_A[0][41] , \cache_data_A[0][40] , \cache_data_A[0][39] ,
         \cache_data_A[0][38] , \cache_data_A[0][37] , \cache_data_A[0][36] ,
         \cache_data_A[0][35] , \cache_data_A[0][34] , \cache_data_A[0][33] ,
         \cache_data_A[0][32] , \cache_data_A[0][31] , \cache_data_A[0][30] ,
         \cache_data_A[0][29] , \cache_data_A[0][28] , \cache_data_A[0][27] ,
         \cache_data_A[0][26] , \cache_data_A[0][25] , \cache_data_A[0][24] ,
         \cache_data_A[0][23] , \cache_data_A[0][22] , \cache_data_A[0][21] ,
         \cache_data_A[0][20] , \cache_data_A[0][19] , \cache_data_A[0][18] ,
         \cache_data_A[0][17] , \cache_data_A[0][16] , \cache_data_A[0][15] ,
         \cache_data_A[0][14] , \cache_data_A[0][13] , \cache_data_A[0][12] ,
         \cache_data_A[0][11] , \cache_data_A[0][10] , \cache_data_A[0][9] ,
         \cache_data_A[0][8] , \cache_data_A[0][7] , \cache_data_A[0][6] ,
         \cache_data_A[0][5] , \cache_data_A[0][4] , \cache_data_A[0][3] ,
         \cache_data_A[0][2] , \cache_data_A[0][1] , \cache_data_A[0][0] ,
         SelectWay, \cache_data_B[7][127] , \cache_data_B[7][126] ,
         \cache_data_B[7][125] , \cache_data_B[7][124] ,
         \cache_data_B[7][123] , \cache_data_B[7][122] ,
         \cache_data_B[7][121] , \cache_data_B[7][120] ,
         \cache_data_B[7][119] , \cache_data_B[7][118] ,
         \cache_data_B[7][117] , \cache_data_B[7][116] ,
         \cache_data_B[7][115] , \cache_data_B[7][114] ,
         \cache_data_B[7][113] , \cache_data_B[7][112] ,
         \cache_data_B[7][111] , \cache_data_B[7][110] ,
         \cache_data_B[7][109] , \cache_data_B[7][108] ,
         \cache_data_B[7][107] , \cache_data_B[7][106] ,
         \cache_data_B[7][105] , \cache_data_B[7][104] ,
         \cache_data_B[7][103] , \cache_data_B[7][102] ,
         \cache_data_B[7][101] , \cache_data_B[7][100] , \cache_data_B[7][99] ,
         \cache_data_B[7][98] , \cache_data_B[7][97] , \cache_data_B[7][96] ,
         \cache_data_B[7][95] , \cache_data_B[7][94] , \cache_data_B[7][93] ,
         \cache_data_B[7][92] , \cache_data_B[7][91] , \cache_data_B[7][90] ,
         \cache_data_B[7][89] , \cache_data_B[7][88] , \cache_data_B[7][87] ,
         \cache_data_B[7][86] , \cache_data_B[7][85] , \cache_data_B[7][84] ,
         \cache_data_B[7][83] , \cache_data_B[7][82] , \cache_data_B[7][81] ,
         \cache_data_B[7][80] , \cache_data_B[7][79] , \cache_data_B[7][78] ,
         \cache_data_B[7][77] , \cache_data_B[7][76] , \cache_data_B[7][75] ,
         \cache_data_B[7][74] , \cache_data_B[7][73] , \cache_data_B[7][72] ,
         \cache_data_B[7][71] , \cache_data_B[7][70] , \cache_data_B[7][69] ,
         \cache_data_B[7][68] , \cache_data_B[7][67] , \cache_data_B[7][66] ,
         \cache_data_B[7][65] , \cache_data_B[7][64] , \cache_data_B[7][63] ,
         \cache_data_B[7][62] , \cache_data_B[7][61] , \cache_data_B[7][60] ,
         \cache_data_B[7][59] , \cache_data_B[7][58] , \cache_data_B[7][57] ,
         \cache_data_B[7][56] , \cache_data_B[7][55] , \cache_data_B[7][54] ,
         \cache_data_B[7][53] , \cache_data_B[7][52] , \cache_data_B[7][51] ,
         \cache_data_B[7][50] , \cache_data_B[7][49] , \cache_data_B[7][48] ,
         \cache_data_B[7][47] , \cache_data_B[7][46] , \cache_data_B[7][45] ,
         \cache_data_B[7][44] , \cache_data_B[7][43] , \cache_data_B[7][42] ,
         \cache_data_B[7][41] , \cache_data_B[7][40] , \cache_data_B[7][39] ,
         \cache_data_B[7][38] , \cache_data_B[7][37] , \cache_data_B[7][36] ,
         \cache_data_B[7][35] , \cache_data_B[7][34] , \cache_data_B[7][33] ,
         \cache_data_B[7][32] , \cache_data_B[7][31] , \cache_data_B[7][30] ,
         \cache_data_B[7][29] , \cache_data_B[7][28] , \cache_data_B[7][27] ,
         \cache_data_B[7][26] , \cache_data_B[7][25] , \cache_data_B[7][24] ,
         \cache_data_B[7][23] , \cache_data_B[7][22] , \cache_data_B[7][21] ,
         \cache_data_B[7][20] , \cache_data_B[7][19] , \cache_data_B[7][18] ,
         \cache_data_B[7][17] , \cache_data_B[7][16] , \cache_data_B[7][15] ,
         \cache_data_B[7][14] , \cache_data_B[7][13] , \cache_data_B[7][12] ,
         \cache_data_B[7][11] , \cache_data_B[7][10] , \cache_data_B[7][9] ,
         \cache_data_B[7][8] , \cache_data_B[7][7] , \cache_data_B[7][6] ,
         \cache_data_B[7][5] , \cache_data_B[7][4] , \cache_data_B[7][3] ,
         \cache_data_B[7][2] , \cache_data_B[7][1] , \cache_data_B[7][0] ,
         \cache_data_B[6][127] , \cache_data_B[6][126] ,
         \cache_data_B[6][125] , \cache_data_B[6][124] ,
         \cache_data_B[6][123] , \cache_data_B[6][122] ,
         \cache_data_B[6][121] , \cache_data_B[6][120] ,
         \cache_data_B[6][119] , \cache_data_B[6][118] ,
         \cache_data_B[6][117] , \cache_data_B[6][116] ,
         \cache_data_B[6][115] , \cache_data_B[6][114] ,
         \cache_data_B[6][113] , \cache_data_B[6][112] ,
         \cache_data_B[6][111] , \cache_data_B[6][110] ,
         \cache_data_B[6][109] , \cache_data_B[6][108] ,
         \cache_data_B[6][107] , \cache_data_B[6][106] ,
         \cache_data_B[6][105] , \cache_data_B[6][104] ,
         \cache_data_B[6][103] , \cache_data_B[6][102] ,
         \cache_data_B[6][101] , \cache_data_B[6][100] , \cache_data_B[6][99] ,
         \cache_data_B[6][98] , \cache_data_B[6][97] , \cache_data_B[6][96] ,
         \cache_data_B[6][95] , \cache_data_B[6][94] , \cache_data_B[6][93] ,
         \cache_data_B[6][92] , \cache_data_B[6][91] , \cache_data_B[6][90] ,
         \cache_data_B[6][89] , \cache_data_B[6][88] , \cache_data_B[6][87] ,
         \cache_data_B[6][86] , \cache_data_B[6][85] , \cache_data_B[6][84] ,
         \cache_data_B[6][83] , \cache_data_B[6][82] , \cache_data_B[6][81] ,
         \cache_data_B[6][80] , \cache_data_B[6][79] , \cache_data_B[6][78] ,
         \cache_data_B[6][77] , \cache_data_B[6][76] , \cache_data_B[6][75] ,
         \cache_data_B[6][74] , \cache_data_B[6][73] , \cache_data_B[6][72] ,
         \cache_data_B[6][71] , \cache_data_B[6][70] , \cache_data_B[6][69] ,
         \cache_data_B[6][68] , \cache_data_B[6][67] , \cache_data_B[6][66] ,
         \cache_data_B[6][65] , \cache_data_B[6][64] , \cache_data_B[6][63] ,
         \cache_data_B[6][62] , \cache_data_B[6][61] , \cache_data_B[6][60] ,
         \cache_data_B[6][59] , \cache_data_B[6][58] , \cache_data_B[6][57] ,
         \cache_data_B[6][56] , \cache_data_B[6][55] , \cache_data_B[6][54] ,
         \cache_data_B[6][53] , \cache_data_B[6][52] , \cache_data_B[6][51] ,
         \cache_data_B[6][50] , \cache_data_B[6][49] , \cache_data_B[6][48] ,
         \cache_data_B[6][47] , \cache_data_B[6][46] , \cache_data_B[6][45] ,
         \cache_data_B[6][44] , \cache_data_B[6][43] , \cache_data_B[6][42] ,
         \cache_data_B[6][41] , \cache_data_B[6][40] , \cache_data_B[6][39] ,
         \cache_data_B[6][38] , \cache_data_B[6][37] , \cache_data_B[6][36] ,
         \cache_data_B[6][35] , \cache_data_B[6][34] , \cache_data_B[6][33] ,
         \cache_data_B[6][32] , \cache_data_B[6][31] , \cache_data_B[6][30] ,
         \cache_data_B[6][29] , \cache_data_B[6][28] , \cache_data_B[6][27] ,
         \cache_data_B[6][26] , \cache_data_B[6][25] , \cache_data_B[6][24] ,
         \cache_data_B[6][23] , \cache_data_B[6][22] , \cache_data_B[6][21] ,
         \cache_data_B[6][20] , \cache_data_B[6][19] , \cache_data_B[6][18] ,
         \cache_data_B[6][17] , \cache_data_B[6][16] , \cache_data_B[6][15] ,
         \cache_data_B[6][14] , \cache_data_B[6][13] , \cache_data_B[6][12] ,
         \cache_data_B[6][11] , \cache_data_B[6][10] , \cache_data_B[6][9] ,
         \cache_data_B[6][8] , \cache_data_B[6][7] , \cache_data_B[6][6] ,
         \cache_data_B[6][5] , \cache_data_B[6][4] , \cache_data_B[6][3] ,
         \cache_data_B[6][2] , \cache_data_B[6][1] , \cache_data_B[6][0] ,
         \cache_data_B[5][127] , \cache_data_B[5][126] ,
         \cache_data_B[5][125] , \cache_data_B[5][124] ,
         \cache_data_B[5][123] , \cache_data_B[5][122] ,
         \cache_data_B[5][121] , \cache_data_B[5][120] ,
         \cache_data_B[5][119] , \cache_data_B[5][118] ,
         \cache_data_B[5][117] , \cache_data_B[5][116] ,
         \cache_data_B[5][115] , \cache_data_B[5][114] ,
         \cache_data_B[5][113] , \cache_data_B[5][112] ,
         \cache_data_B[5][111] , \cache_data_B[5][110] ,
         \cache_data_B[5][109] , \cache_data_B[5][108] ,
         \cache_data_B[5][107] , \cache_data_B[5][106] ,
         \cache_data_B[5][105] , \cache_data_B[5][104] ,
         \cache_data_B[5][103] , \cache_data_B[5][102] ,
         \cache_data_B[5][101] , \cache_data_B[5][100] , \cache_data_B[5][99] ,
         \cache_data_B[5][98] , \cache_data_B[5][97] , \cache_data_B[5][96] ,
         \cache_data_B[5][95] , \cache_data_B[5][94] , \cache_data_B[5][93] ,
         \cache_data_B[5][92] , \cache_data_B[5][91] , \cache_data_B[5][90] ,
         \cache_data_B[5][89] , \cache_data_B[5][88] , \cache_data_B[5][87] ,
         \cache_data_B[5][86] , \cache_data_B[5][85] , \cache_data_B[5][84] ,
         \cache_data_B[5][83] , \cache_data_B[5][82] , \cache_data_B[5][81] ,
         \cache_data_B[5][80] , \cache_data_B[5][79] , \cache_data_B[5][78] ,
         \cache_data_B[5][77] , \cache_data_B[5][76] , \cache_data_B[5][75] ,
         \cache_data_B[5][74] , \cache_data_B[5][73] , \cache_data_B[5][72] ,
         \cache_data_B[5][71] , \cache_data_B[5][70] , \cache_data_B[5][69] ,
         \cache_data_B[5][68] , \cache_data_B[5][67] , \cache_data_B[5][66] ,
         \cache_data_B[5][65] , \cache_data_B[5][64] , \cache_data_B[5][63] ,
         \cache_data_B[5][62] , \cache_data_B[5][61] , \cache_data_B[5][60] ,
         \cache_data_B[5][59] , \cache_data_B[5][58] , \cache_data_B[5][57] ,
         \cache_data_B[5][56] , \cache_data_B[5][55] , \cache_data_B[5][54] ,
         \cache_data_B[5][53] , \cache_data_B[5][52] , \cache_data_B[5][51] ,
         \cache_data_B[5][50] , \cache_data_B[5][49] , \cache_data_B[5][48] ,
         \cache_data_B[5][47] , \cache_data_B[5][46] , \cache_data_B[5][45] ,
         \cache_data_B[5][44] , \cache_data_B[5][43] , \cache_data_B[5][42] ,
         \cache_data_B[5][41] , \cache_data_B[5][40] , \cache_data_B[5][39] ,
         \cache_data_B[5][38] , \cache_data_B[5][37] , \cache_data_B[5][36] ,
         \cache_data_B[5][35] , \cache_data_B[5][34] , \cache_data_B[5][33] ,
         \cache_data_B[5][32] , \cache_data_B[5][31] , \cache_data_B[5][30] ,
         \cache_data_B[5][29] , \cache_data_B[5][28] , \cache_data_B[5][27] ,
         \cache_data_B[5][26] , \cache_data_B[5][25] , \cache_data_B[5][24] ,
         \cache_data_B[5][23] , \cache_data_B[5][22] , \cache_data_B[5][21] ,
         \cache_data_B[5][20] , \cache_data_B[5][19] , \cache_data_B[5][18] ,
         \cache_data_B[5][17] , \cache_data_B[5][16] , \cache_data_B[5][15] ,
         \cache_data_B[5][14] , \cache_data_B[5][13] , \cache_data_B[5][12] ,
         \cache_data_B[5][11] , \cache_data_B[5][10] , \cache_data_B[5][9] ,
         \cache_data_B[5][8] , \cache_data_B[5][7] , \cache_data_B[5][6] ,
         \cache_data_B[5][5] , \cache_data_B[5][4] , \cache_data_B[5][3] ,
         \cache_data_B[5][2] , \cache_data_B[5][1] , \cache_data_B[5][0] ,
         \cache_data_B[4][127] , \cache_data_B[4][126] ,
         \cache_data_B[4][125] , \cache_data_B[4][124] ,
         \cache_data_B[4][123] , \cache_data_B[4][122] ,
         \cache_data_B[4][121] , \cache_data_B[4][120] ,
         \cache_data_B[4][119] , \cache_data_B[4][118] ,
         \cache_data_B[4][117] , \cache_data_B[4][116] ,
         \cache_data_B[4][115] , \cache_data_B[4][114] ,
         \cache_data_B[4][113] , \cache_data_B[4][112] ,
         \cache_data_B[4][111] , \cache_data_B[4][110] ,
         \cache_data_B[4][109] , \cache_data_B[4][108] ,
         \cache_data_B[4][107] , \cache_data_B[4][106] ,
         \cache_data_B[4][105] , \cache_data_B[4][104] ,
         \cache_data_B[4][103] , \cache_data_B[4][102] ,
         \cache_data_B[4][101] , \cache_data_B[4][100] , \cache_data_B[4][99] ,
         \cache_data_B[4][98] , \cache_data_B[4][97] , \cache_data_B[4][96] ,
         \cache_data_B[4][95] , \cache_data_B[4][94] , \cache_data_B[4][93] ,
         \cache_data_B[4][92] , \cache_data_B[4][91] , \cache_data_B[4][90] ,
         \cache_data_B[4][89] , \cache_data_B[4][88] , \cache_data_B[4][87] ,
         \cache_data_B[4][86] , \cache_data_B[4][85] , \cache_data_B[4][84] ,
         \cache_data_B[4][83] , \cache_data_B[4][82] , \cache_data_B[4][81] ,
         \cache_data_B[4][80] , \cache_data_B[4][79] , \cache_data_B[4][78] ,
         \cache_data_B[4][77] , \cache_data_B[4][76] , \cache_data_B[4][75] ,
         \cache_data_B[4][74] , \cache_data_B[4][73] , \cache_data_B[4][72] ,
         \cache_data_B[4][71] , \cache_data_B[4][70] , \cache_data_B[4][69] ,
         \cache_data_B[4][68] , \cache_data_B[4][67] , \cache_data_B[4][66] ,
         \cache_data_B[4][65] , \cache_data_B[4][64] , \cache_data_B[4][63] ,
         \cache_data_B[4][62] , \cache_data_B[4][61] , \cache_data_B[4][60] ,
         \cache_data_B[4][59] , \cache_data_B[4][58] , \cache_data_B[4][57] ,
         \cache_data_B[4][56] , \cache_data_B[4][55] , \cache_data_B[4][54] ,
         \cache_data_B[4][53] , \cache_data_B[4][52] , \cache_data_B[4][51] ,
         \cache_data_B[4][50] , \cache_data_B[4][49] , \cache_data_B[4][48] ,
         \cache_data_B[4][47] , \cache_data_B[4][46] , \cache_data_B[4][45] ,
         \cache_data_B[4][44] , \cache_data_B[4][43] , \cache_data_B[4][42] ,
         \cache_data_B[4][41] , \cache_data_B[4][40] , \cache_data_B[4][39] ,
         \cache_data_B[4][38] , \cache_data_B[4][37] , \cache_data_B[4][36] ,
         \cache_data_B[4][35] , \cache_data_B[4][34] , \cache_data_B[4][33] ,
         \cache_data_B[4][32] , \cache_data_B[4][31] , \cache_data_B[4][30] ,
         \cache_data_B[4][29] , \cache_data_B[4][28] , \cache_data_B[4][27] ,
         \cache_data_B[4][26] , \cache_data_B[4][25] , \cache_data_B[4][24] ,
         \cache_data_B[4][23] , \cache_data_B[4][22] , \cache_data_B[4][21] ,
         \cache_data_B[4][20] , \cache_data_B[4][19] , \cache_data_B[4][18] ,
         \cache_data_B[4][17] , \cache_data_B[4][16] , \cache_data_B[4][15] ,
         \cache_data_B[4][14] , \cache_data_B[4][13] , \cache_data_B[4][12] ,
         \cache_data_B[4][11] , \cache_data_B[4][10] , \cache_data_B[4][9] ,
         \cache_data_B[4][8] , \cache_data_B[4][7] , \cache_data_B[4][6] ,
         \cache_data_B[4][5] , \cache_data_B[4][4] , \cache_data_B[4][3] ,
         \cache_data_B[4][2] , \cache_data_B[4][1] , \cache_data_B[4][0] ,
         \cache_data_B[3][127] , \cache_data_B[3][126] ,
         \cache_data_B[3][125] , \cache_data_B[3][124] ,
         \cache_data_B[3][123] , \cache_data_B[3][122] ,
         \cache_data_B[3][121] , \cache_data_B[3][120] ,
         \cache_data_B[3][119] , \cache_data_B[3][118] ,
         \cache_data_B[3][117] , \cache_data_B[3][116] ,
         \cache_data_B[3][115] , \cache_data_B[3][114] ,
         \cache_data_B[3][113] , \cache_data_B[3][112] ,
         \cache_data_B[3][111] , \cache_data_B[3][110] ,
         \cache_data_B[3][109] , \cache_data_B[3][108] ,
         \cache_data_B[3][107] , \cache_data_B[3][106] ,
         \cache_data_B[3][105] , \cache_data_B[3][104] ,
         \cache_data_B[3][103] , \cache_data_B[3][102] ,
         \cache_data_B[3][101] , \cache_data_B[3][100] , \cache_data_B[3][99] ,
         \cache_data_B[3][98] , \cache_data_B[3][97] , \cache_data_B[3][96] ,
         \cache_data_B[3][95] , \cache_data_B[3][94] , \cache_data_B[3][93] ,
         \cache_data_B[3][92] , \cache_data_B[3][91] , \cache_data_B[3][90] ,
         \cache_data_B[3][89] , \cache_data_B[3][88] , \cache_data_B[3][87] ,
         \cache_data_B[3][86] , \cache_data_B[3][85] , \cache_data_B[3][84] ,
         \cache_data_B[3][83] , \cache_data_B[3][82] , \cache_data_B[3][81] ,
         \cache_data_B[3][80] , \cache_data_B[3][79] , \cache_data_B[3][78] ,
         \cache_data_B[3][77] , \cache_data_B[3][76] , \cache_data_B[3][75] ,
         \cache_data_B[3][74] , \cache_data_B[3][73] , \cache_data_B[3][72] ,
         \cache_data_B[3][71] , \cache_data_B[3][70] , \cache_data_B[3][69] ,
         \cache_data_B[3][68] , \cache_data_B[3][67] , \cache_data_B[3][66] ,
         \cache_data_B[3][65] , \cache_data_B[3][64] , \cache_data_B[3][63] ,
         \cache_data_B[3][62] , \cache_data_B[3][61] , \cache_data_B[3][60] ,
         \cache_data_B[3][59] , \cache_data_B[3][58] , \cache_data_B[3][57] ,
         \cache_data_B[3][56] , \cache_data_B[3][55] , \cache_data_B[3][54] ,
         \cache_data_B[3][53] , \cache_data_B[3][52] , \cache_data_B[3][51] ,
         \cache_data_B[3][50] , \cache_data_B[3][49] , \cache_data_B[3][48] ,
         \cache_data_B[3][47] , \cache_data_B[3][46] , \cache_data_B[3][45] ,
         \cache_data_B[3][44] , \cache_data_B[3][43] , \cache_data_B[3][42] ,
         \cache_data_B[3][41] , \cache_data_B[3][40] , \cache_data_B[3][39] ,
         \cache_data_B[3][38] , \cache_data_B[3][37] , \cache_data_B[3][36] ,
         \cache_data_B[3][35] , \cache_data_B[3][34] , \cache_data_B[3][33] ,
         \cache_data_B[3][32] , \cache_data_B[3][31] , \cache_data_B[3][30] ,
         \cache_data_B[3][29] , \cache_data_B[3][28] , \cache_data_B[3][27] ,
         \cache_data_B[3][26] , \cache_data_B[3][25] , \cache_data_B[3][24] ,
         \cache_data_B[3][23] , \cache_data_B[3][22] , \cache_data_B[3][21] ,
         \cache_data_B[3][20] , \cache_data_B[3][19] , \cache_data_B[3][18] ,
         \cache_data_B[3][17] , \cache_data_B[3][16] , \cache_data_B[3][15] ,
         \cache_data_B[3][14] , \cache_data_B[3][13] , \cache_data_B[3][12] ,
         \cache_data_B[3][11] , \cache_data_B[3][10] , \cache_data_B[3][9] ,
         \cache_data_B[3][8] , \cache_data_B[3][7] , \cache_data_B[3][6] ,
         \cache_data_B[3][5] , \cache_data_B[3][4] , \cache_data_B[3][3] ,
         \cache_data_B[3][2] , \cache_data_B[3][1] , \cache_data_B[3][0] ,
         \cache_data_B[2][127] , \cache_data_B[2][126] ,
         \cache_data_B[2][125] , \cache_data_B[2][124] ,
         \cache_data_B[2][123] , \cache_data_B[2][122] ,
         \cache_data_B[2][121] , \cache_data_B[2][120] ,
         \cache_data_B[2][119] , \cache_data_B[2][118] ,
         \cache_data_B[2][117] , \cache_data_B[2][116] ,
         \cache_data_B[2][115] , \cache_data_B[2][114] ,
         \cache_data_B[2][113] , \cache_data_B[2][112] ,
         \cache_data_B[2][111] , \cache_data_B[2][110] ,
         \cache_data_B[2][109] , \cache_data_B[2][108] ,
         \cache_data_B[2][107] , \cache_data_B[2][106] ,
         \cache_data_B[2][105] , \cache_data_B[2][104] ,
         \cache_data_B[2][103] , \cache_data_B[2][102] ,
         \cache_data_B[2][101] , \cache_data_B[2][100] , \cache_data_B[2][99] ,
         \cache_data_B[2][98] , \cache_data_B[2][97] , \cache_data_B[2][96] ,
         \cache_data_B[2][95] , \cache_data_B[2][94] , \cache_data_B[2][93] ,
         \cache_data_B[2][92] , \cache_data_B[2][91] , \cache_data_B[2][90] ,
         \cache_data_B[2][89] , \cache_data_B[2][88] , \cache_data_B[2][87] ,
         \cache_data_B[2][86] , \cache_data_B[2][85] , \cache_data_B[2][84] ,
         \cache_data_B[2][83] , \cache_data_B[2][82] , \cache_data_B[2][81] ,
         \cache_data_B[2][80] , \cache_data_B[2][79] , \cache_data_B[2][78] ,
         \cache_data_B[2][77] , \cache_data_B[2][76] , \cache_data_B[2][75] ,
         \cache_data_B[2][74] , \cache_data_B[2][73] , \cache_data_B[2][72] ,
         \cache_data_B[2][71] , \cache_data_B[2][70] , \cache_data_B[2][69] ,
         \cache_data_B[2][68] , \cache_data_B[2][67] , \cache_data_B[2][66] ,
         \cache_data_B[2][65] , \cache_data_B[2][64] , \cache_data_B[2][63] ,
         \cache_data_B[2][62] , \cache_data_B[2][61] , \cache_data_B[2][60] ,
         \cache_data_B[2][59] , \cache_data_B[2][58] , \cache_data_B[2][57] ,
         \cache_data_B[2][56] , \cache_data_B[2][55] , \cache_data_B[2][54] ,
         \cache_data_B[2][53] , \cache_data_B[2][52] , \cache_data_B[2][51] ,
         \cache_data_B[2][50] , \cache_data_B[2][49] , \cache_data_B[2][48] ,
         \cache_data_B[2][47] , \cache_data_B[2][46] , \cache_data_B[2][45] ,
         \cache_data_B[2][44] , \cache_data_B[2][43] , \cache_data_B[2][42] ,
         \cache_data_B[2][41] , \cache_data_B[2][40] , \cache_data_B[2][39] ,
         \cache_data_B[2][38] , \cache_data_B[2][37] , \cache_data_B[2][36] ,
         \cache_data_B[2][35] , \cache_data_B[2][34] , \cache_data_B[2][33] ,
         \cache_data_B[2][32] , \cache_data_B[2][31] , \cache_data_B[2][30] ,
         \cache_data_B[2][29] , \cache_data_B[2][28] , \cache_data_B[2][27] ,
         \cache_data_B[2][26] , \cache_data_B[2][25] , \cache_data_B[2][24] ,
         \cache_data_B[2][23] , \cache_data_B[2][22] , \cache_data_B[2][21] ,
         \cache_data_B[2][20] , \cache_data_B[2][19] , \cache_data_B[2][18] ,
         \cache_data_B[2][17] , \cache_data_B[2][16] , \cache_data_B[2][15] ,
         \cache_data_B[2][14] , \cache_data_B[2][13] , \cache_data_B[2][12] ,
         \cache_data_B[2][11] , \cache_data_B[2][10] , \cache_data_B[2][9] ,
         \cache_data_B[2][8] , \cache_data_B[2][7] , \cache_data_B[2][6] ,
         \cache_data_B[2][5] , \cache_data_B[2][4] , \cache_data_B[2][3] ,
         \cache_data_B[2][2] , \cache_data_B[2][1] , \cache_data_B[2][0] ,
         \cache_data_B[1][127] , \cache_data_B[1][126] ,
         \cache_data_B[1][125] , \cache_data_B[1][124] ,
         \cache_data_B[1][123] , \cache_data_B[1][122] ,
         \cache_data_B[1][121] , \cache_data_B[1][120] ,
         \cache_data_B[1][119] , \cache_data_B[1][118] ,
         \cache_data_B[1][117] , \cache_data_B[1][116] ,
         \cache_data_B[1][115] , \cache_data_B[1][114] ,
         \cache_data_B[1][113] , \cache_data_B[1][112] ,
         \cache_data_B[1][111] , \cache_data_B[1][110] ,
         \cache_data_B[1][109] , \cache_data_B[1][108] ,
         \cache_data_B[1][107] , \cache_data_B[1][106] ,
         \cache_data_B[1][105] , \cache_data_B[1][104] ,
         \cache_data_B[1][103] , \cache_data_B[1][102] ,
         \cache_data_B[1][101] , \cache_data_B[1][100] , \cache_data_B[1][99] ,
         \cache_data_B[1][98] , \cache_data_B[1][97] , \cache_data_B[1][96] ,
         \cache_data_B[1][95] , \cache_data_B[1][94] , \cache_data_B[1][93] ,
         \cache_data_B[1][92] , \cache_data_B[1][91] , \cache_data_B[1][90] ,
         \cache_data_B[1][89] , \cache_data_B[1][88] , \cache_data_B[1][87] ,
         \cache_data_B[1][86] , \cache_data_B[1][85] , \cache_data_B[1][84] ,
         \cache_data_B[1][83] , \cache_data_B[1][82] , \cache_data_B[1][81] ,
         \cache_data_B[1][80] , \cache_data_B[1][79] , \cache_data_B[1][78] ,
         \cache_data_B[1][77] , \cache_data_B[1][76] , \cache_data_B[1][75] ,
         \cache_data_B[1][74] , \cache_data_B[1][73] , \cache_data_B[1][72] ,
         \cache_data_B[1][71] , \cache_data_B[1][70] , \cache_data_B[1][69] ,
         \cache_data_B[1][68] , \cache_data_B[1][67] , \cache_data_B[1][66] ,
         \cache_data_B[1][65] , \cache_data_B[1][64] , \cache_data_B[1][63] ,
         \cache_data_B[1][62] , \cache_data_B[1][61] , \cache_data_B[1][60] ,
         \cache_data_B[1][59] , \cache_data_B[1][58] , \cache_data_B[1][57] ,
         \cache_data_B[1][56] , \cache_data_B[1][55] , \cache_data_B[1][54] ,
         \cache_data_B[1][53] , \cache_data_B[1][52] , \cache_data_B[1][51] ,
         \cache_data_B[1][50] , \cache_data_B[1][49] , \cache_data_B[1][48] ,
         \cache_data_B[1][47] , \cache_data_B[1][46] , \cache_data_B[1][45] ,
         \cache_data_B[1][44] , \cache_data_B[1][43] , \cache_data_B[1][42] ,
         \cache_data_B[1][41] , \cache_data_B[1][40] , \cache_data_B[1][39] ,
         \cache_data_B[1][38] , \cache_data_B[1][37] , \cache_data_B[1][36] ,
         \cache_data_B[1][35] , \cache_data_B[1][34] , \cache_data_B[1][33] ,
         \cache_data_B[1][32] , \cache_data_B[1][31] , \cache_data_B[1][30] ,
         \cache_data_B[1][29] , \cache_data_B[1][28] , \cache_data_B[1][27] ,
         \cache_data_B[1][26] , \cache_data_B[1][25] , \cache_data_B[1][24] ,
         \cache_data_B[1][23] , \cache_data_B[1][22] , \cache_data_B[1][21] ,
         \cache_data_B[1][20] , \cache_data_B[1][19] , \cache_data_B[1][18] ,
         \cache_data_B[1][17] , \cache_data_B[1][16] , \cache_data_B[1][15] ,
         \cache_data_B[1][14] , \cache_data_B[1][13] , \cache_data_B[1][12] ,
         \cache_data_B[1][11] , \cache_data_B[1][10] , \cache_data_B[1][9] ,
         \cache_data_B[1][8] , \cache_data_B[1][7] , \cache_data_B[1][6] ,
         \cache_data_B[1][5] , \cache_data_B[1][4] , \cache_data_B[1][3] ,
         \cache_data_B[1][2] , \cache_data_B[1][1] , \cache_data_B[1][0] ,
         \cache_data_B[0][127] , \cache_data_B[0][126] ,
         \cache_data_B[0][125] , \cache_data_B[0][124] ,
         \cache_data_B[0][123] , \cache_data_B[0][122] ,
         \cache_data_B[0][121] , \cache_data_B[0][120] ,
         \cache_data_B[0][119] , \cache_data_B[0][118] ,
         \cache_data_B[0][117] , \cache_data_B[0][116] ,
         \cache_data_B[0][115] , \cache_data_B[0][114] ,
         \cache_data_B[0][113] , \cache_data_B[0][112] ,
         \cache_data_B[0][111] , \cache_data_B[0][110] ,
         \cache_data_B[0][109] , \cache_data_B[0][108] ,
         \cache_data_B[0][107] , \cache_data_B[0][106] ,
         \cache_data_B[0][105] , \cache_data_B[0][104] ,
         \cache_data_B[0][103] , \cache_data_B[0][102] ,
         \cache_data_B[0][101] , \cache_data_B[0][100] , \cache_data_B[0][99] ,
         \cache_data_B[0][98] , \cache_data_B[0][97] , \cache_data_B[0][96] ,
         \cache_data_B[0][95] , \cache_data_B[0][94] , \cache_data_B[0][93] ,
         \cache_data_B[0][92] , \cache_data_B[0][91] , \cache_data_B[0][90] ,
         \cache_data_B[0][89] , \cache_data_B[0][88] , \cache_data_B[0][87] ,
         \cache_data_B[0][86] , \cache_data_B[0][85] , \cache_data_B[0][84] ,
         \cache_data_B[0][83] , \cache_data_B[0][82] , \cache_data_B[0][81] ,
         \cache_data_B[0][80] , \cache_data_B[0][79] , \cache_data_B[0][78] ,
         \cache_data_B[0][77] , \cache_data_B[0][76] , \cache_data_B[0][75] ,
         \cache_data_B[0][74] , \cache_data_B[0][73] , \cache_data_B[0][72] ,
         \cache_data_B[0][71] , \cache_data_B[0][70] , \cache_data_B[0][69] ,
         \cache_data_B[0][68] , \cache_data_B[0][67] , \cache_data_B[0][66] ,
         \cache_data_B[0][65] , \cache_data_B[0][64] , \cache_data_B[0][63] ,
         \cache_data_B[0][62] , \cache_data_B[0][61] , \cache_data_B[0][60] ,
         \cache_data_B[0][59] , \cache_data_B[0][58] , \cache_data_B[0][57] ,
         \cache_data_B[0][56] , \cache_data_B[0][55] , \cache_data_B[0][54] ,
         \cache_data_B[0][53] , \cache_data_B[0][52] , \cache_data_B[0][51] ,
         \cache_data_B[0][50] , \cache_data_B[0][49] , \cache_data_B[0][48] ,
         \cache_data_B[0][47] , \cache_data_B[0][46] , \cache_data_B[0][45] ,
         \cache_data_B[0][44] , \cache_data_B[0][43] , \cache_data_B[0][42] ,
         \cache_data_B[0][41] , \cache_data_B[0][40] , \cache_data_B[0][39] ,
         \cache_data_B[0][38] , \cache_data_B[0][37] , \cache_data_B[0][36] ,
         \cache_data_B[0][35] , \cache_data_B[0][34] , \cache_data_B[0][33] ,
         \cache_data_B[0][32] , \cache_data_B[0][31] , \cache_data_B[0][30] ,
         \cache_data_B[0][29] , \cache_data_B[0][28] , \cache_data_B[0][27] ,
         \cache_data_B[0][26] , \cache_data_B[0][25] , \cache_data_B[0][24] ,
         \cache_data_B[0][23] , \cache_data_B[0][22] , \cache_data_B[0][21] ,
         \cache_data_B[0][20] , \cache_data_B[0][19] , \cache_data_B[0][18] ,
         \cache_data_B[0][17] , \cache_data_B[0][16] , \cache_data_B[0][15] ,
         \cache_data_B[0][14] , \cache_data_B[0][13] , \cache_data_B[0][12] ,
         \cache_data_B[0][11] , \cache_data_B[0][10] , \cache_data_B[0][9] ,
         \cache_data_B[0][8] , \cache_data_B[0][7] , \cache_data_B[0][6] ,
         \cache_data_B[0][5] , \cache_data_B[0][4] , \cache_data_B[0][3] ,
         \cache_data_B[0][2] , \cache_data_B[0][1] , \cache_data_B[0][0] ,
         rd_temp, \cache_tag_B[7][24] , \cache_tag_B[7][23] ,
         \cache_tag_B[7][22] , \cache_tag_B[7][21] , \cache_tag_B[7][20] ,
         \cache_tag_B[7][19] , \cache_tag_B[7][18] , \cache_tag_B[7][17] ,
         \cache_tag_B[7][16] , \cache_tag_B[7][15] , \cache_tag_B[7][14] ,
         \cache_tag_B[7][13] , \cache_tag_B[7][12] , \cache_tag_B[7][11] ,
         \cache_tag_B[7][10] , \cache_tag_B[7][9] , \cache_tag_B[7][8] ,
         \cache_tag_B[7][7] , \cache_tag_B[7][6] , \cache_tag_B[7][5] ,
         \cache_tag_B[7][4] , \cache_tag_B[7][3] , \cache_tag_B[7][2] ,
         \cache_tag_B[7][1] , \cache_tag_B[7][0] , \cache_tag_B[6][24] ,
         \cache_tag_B[6][23] , \cache_tag_B[6][22] , \cache_tag_B[6][21] ,
         \cache_tag_B[6][20] , \cache_tag_B[6][19] , \cache_tag_B[6][18] ,
         \cache_tag_B[6][17] , \cache_tag_B[6][16] , \cache_tag_B[6][15] ,
         \cache_tag_B[6][14] , \cache_tag_B[6][13] , \cache_tag_B[6][12] ,
         \cache_tag_B[6][11] , \cache_tag_B[6][10] , \cache_tag_B[6][9] ,
         \cache_tag_B[6][8] , \cache_tag_B[6][7] , \cache_tag_B[6][6] ,
         \cache_tag_B[6][5] , \cache_tag_B[6][4] , \cache_tag_B[6][3] ,
         \cache_tag_B[6][2] , \cache_tag_B[6][1] , \cache_tag_B[6][0] ,
         \cache_tag_B[5][24] , \cache_tag_B[5][23] , \cache_tag_B[5][22] ,
         \cache_tag_B[5][21] , \cache_tag_B[5][20] , \cache_tag_B[5][19] ,
         \cache_tag_B[5][18] , \cache_tag_B[5][17] , \cache_tag_B[5][16] ,
         \cache_tag_B[5][15] , \cache_tag_B[5][14] , \cache_tag_B[5][13] ,
         \cache_tag_B[5][12] , \cache_tag_B[5][11] , \cache_tag_B[5][10] ,
         \cache_tag_B[5][9] , \cache_tag_B[5][8] , \cache_tag_B[5][7] ,
         \cache_tag_B[5][6] , \cache_tag_B[5][5] , \cache_tag_B[5][4] ,
         \cache_tag_B[5][3] , \cache_tag_B[5][2] , \cache_tag_B[5][1] ,
         \cache_tag_B[5][0] , \cache_tag_B[4][24] , \cache_tag_B[4][23] ,
         \cache_tag_B[4][22] , \cache_tag_B[4][21] , \cache_tag_B[4][20] ,
         \cache_tag_B[4][19] , \cache_tag_B[4][18] , \cache_tag_B[4][17] ,
         \cache_tag_B[4][16] , \cache_tag_B[4][15] , \cache_tag_B[4][14] ,
         \cache_tag_B[4][13] , \cache_tag_B[4][12] , \cache_tag_B[4][11] ,
         \cache_tag_B[4][10] , \cache_tag_B[4][9] , \cache_tag_B[4][8] ,
         \cache_tag_B[4][7] , \cache_tag_B[4][6] , \cache_tag_B[4][5] ,
         \cache_tag_B[4][4] , \cache_tag_B[4][3] , \cache_tag_B[4][2] ,
         \cache_tag_B[4][1] , \cache_tag_B[4][0] , \cache_tag_B[3][24] ,
         \cache_tag_B[3][23] , \cache_tag_B[3][22] , \cache_tag_B[3][21] ,
         \cache_tag_B[3][20] , \cache_tag_B[3][19] , \cache_tag_B[3][18] ,
         \cache_tag_B[3][17] , \cache_tag_B[3][16] , \cache_tag_B[3][15] ,
         \cache_tag_B[3][14] , \cache_tag_B[3][13] , \cache_tag_B[3][12] ,
         \cache_tag_B[3][11] , \cache_tag_B[3][10] , \cache_tag_B[3][9] ,
         \cache_tag_B[3][8] , \cache_tag_B[3][7] , \cache_tag_B[3][6] ,
         \cache_tag_B[3][5] , \cache_tag_B[3][4] , \cache_tag_B[3][3] ,
         \cache_tag_B[3][2] , \cache_tag_B[3][1] , \cache_tag_B[3][0] ,
         \cache_tag_B[2][24] , \cache_tag_B[2][23] , \cache_tag_B[2][22] ,
         \cache_tag_B[2][21] , \cache_tag_B[2][20] , \cache_tag_B[2][19] ,
         \cache_tag_B[2][18] , \cache_tag_B[2][17] , \cache_tag_B[2][16] ,
         \cache_tag_B[2][15] , \cache_tag_B[2][14] , \cache_tag_B[2][13] ,
         \cache_tag_B[2][12] , \cache_tag_B[2][11] , \cache_tag_B[2][10] ,
         \cache_tag_B[2][9] , \cache_tag_B[2][8] , \cache_tag_B[2][7] ,
         \cache_tag_B[2][6] , \cache_tag_B[2][5] , \cache_tag_B[2][4] ,
         \cache_tag_B[2][3] , \cache_tag_B[2][2] , \cache_tag_B[2][1] ,
         \cache_tag_B[2][0] , \cache_tag_B[1][24] , \cache_tag_B[1][23] ,
         \cache_tag_B[1][22] , \cache_tag_B[1][21] , \cache_tag_B[1][20] ,
         \cache_tag_B[1][19] , \cache_tag_B[1][18] , \cache_tag_B[1][17] ,
         \cache_tag_B[1][16] , \cache_tag_B[1][15] , \cache_tag_B[1][14] ,
         \cache_tag_B[1][13] , \cache_tag_B[1][12] , \cache_tag_B[1][11] ,
         \cache_tag_B[1][10] , \cache_tag_B[1][9] , \cache_tag_B[1][8] ,
         \cache_tag_B[1][7] , \cache_tag_B[1][6] , \cache_tag_B[1][5] ,
         \cache_tag_B[1][4] , \cache_tag_B[1][3] , \cache_tag_B[1][2] ,
         \cache_tag_B[1][1] , \cache_tag_B[1][0] , \cache_tag_B[0][24] ,
         \cache_tag_B[0][23] , \cache_tag_B[0][22] , \cache_tag_B[0][21] ,
         \cache_tag_B[0][20] , \cache_tag_B[0][19] , \cache_tag_B[0][18] ,
         \cache_tag_B[0][17] , \cache_tag_B[0][16] , \cache_tag_B[0][15] ,
         \cache_tag_B[0][14] , \cache_tag_B[0][13] , \cache_tag_B[0][12] ,
         \cache_tag_B[0][11] , \cache_tag_B[0][10] , \cache_tag_B[0][9] ,
         \cache_tag_B[0][8] , \cache_tag_B[0][7] , \cache_tag_B[0][6] ,
         \cache_tag_B[0][5] , \cache_tag_B[0][4] , \cache_tag_B[0][3] ,
         \cache_tag_B[0][2] , \cache_tag_B[0][1] , \cache_tag_B[0][0] , N4111,
         N4112, N4114, N4115, N4117, N4118, N4120, N4121, N4123, N4124, N4126,
         N4127, N4129, N4130, N4132, N4133, N4135, N4136, N4138, N4139, N4141,
         N4142, N4144, N4145, N4147, N4148, N4150, N4151, N4153, N4154, N4156,
         N4157, N4159, N4160, N4162, N4163, N4165, N4166, N4168, N4169, N4171,
         N4172, N4174, N4175, N4177, N4178, N4180, N4181, N4183, N4184, N4186,
         N4187, N4189, N4190, N4192, N4193, N4195, N4196, N4198, N4199, N4201,
         N4202, N4204, N4205, N4207, N4208, N4210, N4211, N4213, N4214, N4216,
         N4217, N4219, N4220, N4222, N4223, N4225, N4226, N4228, N4229, N4231,
         N4232, N4234, N4235, N4237, N4238, N4240, N4241, N4243, N4244, N4246,
         N4247, N4249, N4250, N4252, N4253, N4255, N4256, N4258, N4259, N4261,
         N4262, N4264, N4265, N4267, N4268, N4270, N4271, N4273, N4274, N4276,
         N4277, N4279, N4280, N4282, N4283, N4285, N4286, N4288, N4289, N4291,
         N4292, N4294, N4295, N4297, N4298, N4300, N4301, N4447, N4454, n1, n3,
         n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59,
         n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87,
         n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111,
         n113, n115, n117, n119, n121, n123, n125, n127, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13293, n13294, n13295, n13296, n13297,
         n13298;
  wire   [4:0] state;
  wire   [4:0] next_state;
  wire   [3:0] mem_data_cnt;
  wire   [31:0] iCache_data_wr;
  wire   [7:0] cache_dirty_A;
  wire   [7:0] cache_dirty_B;
  wire   [7:0] cache_valid_A;
  wire   [7:0] cache_valid_B;
  wire   [7:0] cache_line_count;
  assign addr_mem[0] = 1'b0;
  assign addr_mem[1] = 1'b0;

  drsp_1 mem_done_reg ( .ip(N4454), .ck(clk), .rb(1'b1), .s(rst), .q(mem_done)
         );
  drsp_1 \state_reg[0]  ( .ip(next_state[0]), .ck(clk), .rb(1'b1), .s(rst), 
        .q(state[0]) );
  drsp_1 rd_temp_reg ( .ip(n7939), .ck(clk), .rb(1'b1), .s(n13296), .q(rd_temp) );
  drsp_1 \addr_resp_tri_enable_reg[0]  ( .ip(n7937), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4301) );
  drsp_1 \addr_resp_tri_enable_reg[1]  ( .ip(n7935), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4298) );
  drsp_1 \addr_resp_tri_enable_reg[2]  ( .ip(n7933), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4295) );
  drsp_1 \addr_resp_tri_enable_reg[3]  ( .ip(n7931), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4292) );
  drsp_1 \addr_resp_tri_enable_reg[4]  ( .ip(n7929), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4289) );
  drsp_1 \addr_resp_tri_enable_reg[5]  ( .ip(n7927), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4286) );
  drsp_1 \addr_resp_tri_enable_reg[6]  ( .ip(n7925), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4283) );
  drsp_1 \addr_resp_tri_enable_reg[7]  ( .ip(n7899), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4280) );
  drsp_1 \addr_resp_tri_enable_reg[8]  ( .ip(n7881), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4277) );
  drsp_1 \addr_resp_tri_enable_reg[9]  ( .ip(n7863), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4274) );
  drsp_1 \addr_resp_tri_enable_reg[10]  ( .ip(n7845), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4271) );
  drsp_1 \addr_resp_tri_enable_reg[11]  ( .ip(n7827), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4268) );
  drsp_1 \addr_resp_tri_enable_reg[12]  ( .ip(n7809), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4265) );
  drsp_1 \addr_resp_tri_enable_reg[13]  ( .ip(n7791), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4262) );
  drsp_1 \addr_resp_tri_enable_reg[14]  ( .ip(n7773), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4259) );
  drsp_1 \addr_resp_tri_enable_reg[15]  ( .ip(n7755), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4256) );
  drsp_1 \addr_resp_tri_enable_reg[16]  ( .ip(n7737), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4253) );
  drsp_1 \addr_resp_tri_enable_reg[17]  ( .ip(n7719), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4250) );
  drsp_1 \addr_resp_tri_enable_reg[18]  ( .ip(n7701), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4247) );
  drsp_1 \addr_resp_tri_enable_reg[19]  ( .ip(n7683), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4244) );
  drsp_1 \addr_resp_tri_enable_reg[20]  ( .ip(n7665), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4241) );
  drsp_1 \addr_resp_tri_enable_reg[21]  ( .ip(n7647), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4238) );
  drsp_1 \addr_resp_tri_enable_reg[22]  ( .ip(n7629), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4235) );
  drsp_1 \addr_resp_tri_enable_reg[23]  ( .ip(n7611), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4232) );
  drsp_1 \addr_resp_tri_enable_reg[24]  ( .ip(n7593), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4229) );
  drsp_1 \addr_resp_tri_enable_reg[25]  ( .ip(n7575), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4226) );
  drsp_1 \addr_resp_tri_enable_reg[26]  ( .ip(n7557), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4223) );
  drsp_1 \addr_resp_tri_enable_reg[27]  ( .ip(n7539), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4220) );
  drsp_1 \addr_resp_tri_enable_reg[28]  ( .ip(n7521), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4217) );
  drsp_1 \addr_resp_tri_enable_reg[29]  ( .ip(n7503), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4214) );
  drsp_1 \addr_resp_tri_enable_reg[30]  ( .ip(n7485), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4211) );
  drsp_1 \addr_resp_tri_enable_reg[31]  ( .ip(n7467), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4208) );
  drsp_1 busy_reg ( .ip(N4447), .ck(clk), .rb(1'b1), .s(n13298), .q(busy) );
  drsp_1 \data_rd_tri_enable_reg[0]  ( .ip(n7418), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4205) );
  drsp_1 \data_rd_tri_enable_reg[1]  ( .ip(n7417), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4202) );
  drsp_1 \data_rd_tri_enable_reg[2]  ( .ip(n7416), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4199) );
  drsp_1 \data_rd_tri_enable_reg[3]  ( .ip(n7415), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4196) );
  drsp_1 \data_rd_tri_enable_reg[4]  ( .ip(n7414), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4193) );
  drsp_1 \data_rd_tri_enable_reg[5]  ( .ip(n7413), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4190) );
  drsp_1 \data_rd_tri_enable_reg[6]  ( .ip(n7412), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4187) );
  drsp_1 \data_rd_tri_enable_reg[7]  ( .ip(n7411), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4184) );
  drsp_1 \data_rd_tri_enable_reg[8]  ( .ip(n7410), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4181) );
  drsp_1 \data_rd_tri_enable_reg[9]  ( .ip(n7409), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4178) );
  drsp_1 \data_rd_tri_enable_reg[10]  ( .ip(n7408), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4175) );
  drsp_1 \data_rd_tri_enable_reg[11]  ( .ip(n7407), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4172) );
  drsp_1 \data_rd_tri_enable_reg[12]  ( .ip(n7406), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4169) );
  drsp_1 \data_rd_tri_enable_reg[13]  ( .ip(n7405), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4166) );
  drsp_1 \data_rd_tri_enable_reg[14]  ( .ip(n7404), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4163) );
  drsp_1 \data_rd_tri_enable_reg[15]  ( .ip(n7403), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4160) );
  drsp_1 \data_rd_tri_enable_reg[16]  ( .ip(n7402), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4157) );
  drsp_1 \data_rd_tri_enable_reg[17]  ( .ip(n7401), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4154) );
  drsp_1 \data_rd_tri_enable_reg[18]  ( .ip(n7400), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4151) );
  drsp_1 \data_rd_tri_enable_reg[19]  ( .ip(n7399), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4148) );
  drsp_1 \data_rd_tri_enable_reg[20]  ( .ip(n7398), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4145) );
  drsp_1 \data_rd_tri_enable_reg[21]  ( .ip(n7397), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4142) );
  drsp_1 \data_rd_tri_enable_reg[22]  ( .ip(n7396), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4139) );
  drsp_1 \data_rd_tri_enable_reg[23]  ( .ip(n7395), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4136) );
  drsp_1 \data_rd_tri_enable_reg[24]  ( .ip(n7394), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4133) );
  drsp_1 \data_rd_tri_enable_reg[25]  ( .ip(n7393), .ck(clk), .rb(1'b1), .s(
        n13298), .q(N4130) );
  drsp_1 \data_rd_tri_enable_reg[26]  ( .ip(n7392), .ck(clk), .rb(1'b1), .s(
        n13297), .q(N4127) );
  drsp_1 \data_rd_tri_enable_reg[27]  ( .ip(n7391), .ck(clk), .rb(1'b1), .s(
        n13296), .q(N4124) );
  drsp_1 \data_rd_tri_enable_reg[28]  ( .ip(n7390), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4121) );
  drsp_1 \data_rd_tri_enable_reg[29]  ( .ip(n7389), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4118) );
  drsp_1 \data_rd_tri_enable_reg[30]  ( .ip(n7388), .ck(clk), .rb(1'b1), .s(
        n12618), .q(N4115) );
  drsp_1 \data_rd_tri_enable_reg[31]  ( .ip(n7387), .ck(clk), .rb(1'b1), .s(
        rst), .q(N4112) );
  dp_1 SelectWay_reg ( .ip(n7940), .ck(clk), .q(SelectWay) );
  dp_1 \addr_resp_reg[0]  ( .ip(n7938), .ck(clk), .q(N4300) );
  dp_1 \addr_resp_reg[1]  ( .ip(n7936), .ck(clk), .q(N4297) );
  dp_1 \addr_resp_reg[2]  ( .ip(n7934), .ck(clk), .q(N4294) );
  dp_1 \addr_resp_reg[3]  ( .ip(n7932), .ck(clk), .q(N4291) );
  dp_1 \addr_resp_reg[4]  ( .ip(n7930), .ck(clk), .q(N4288) );
  dp_1 \addr_resp_reg[5]  ( .ip(n7928), .ck(clk), .q(N4285) );
  dp_1 \addr_resp_reg[6]  ( .ip(n7926), .ck(clk), .q(N4282) );
  dp_1 \addr_resp_reg[7]  ( .ip(n7900), .ck(clk), .q(N4279) );
  dp_1 \addr_resp_reg[8]  ( .ip(n7882), .ck(clk), .q(N4276) );
  dp_1 \addr_resp_reg[9]  ( .ip(n7864), .ck(clk), .q(N4273) );
  dp_1 \addr_resp_reg[10]  ( .ip(n7846), .ck(clk), .q(N4270) );
  dp_1 \addr_resp_reg[11]  ( .ip(n7828), .ck(clk), .q(N4267) );
  dp_1 \addr_resp_reg[12]  ( .ip(n7810), .ck(clk), .q(N4264) );
  dp_1 \addr_resp_reg[13]  ( .ip(n7792), .ck(clk), .q(N4261) );
  dp_1 \addr_resp_reg[14]  ( .ip(n7774), .ck(clk), .q(N4258) );
  dp_1 \addr_resp_reg[15]  ( .ip(n7756), .ck(clk), .q(N4255) );
  dp_1 \addr_resp_reg[16]  ( .ip(n7738), .ck(clk), .q(N4252) );
  dp_1 \addr_resp_reg[17]  ( .ip(n7720), .ck(clk), .q(N4249) );
  dp_1 \addr_resp_reg[18]  ( .ip(n7702), .ck(clk), .q(N4246) );
  dp_1 \addr_resp_reg[19]  ( .ip(n7684), .ck(clk), .q(N4243) );
  dp_1 \addr_resp_reg[20]  ( .ip(n7666), .ck(clk), .q(N4240) );
  dp_1 \addr_resp_reg[21]  ( .ip(n7648), .ck(clk), .q(N4237) );
  dp_1 \addr_resp_reg[22]  ( .ip(n7630), .ck(clk), .q(N4234) );
  dp_1 \addr_resp_reg[23]  ( .ip(n7612), .ck(clk), .q(N4231) );
  dp_1 \addr_resp_reg[24]  ( .ip(n7594), .ck(clk), .q(N4228) );
  dp_1 \addr_resp_reg[25]  ( .ip(n7576), .ck(clk), .q(N4225) );
  dp_1 \addr_resp_reg[26]  ( .ip(n7558), .ck(clk), .q(N4222) );
  dp_1 \addr_resp_reg[27]  ( .ip(n7540), .ck(clk), .q(N4219) );
  dp_1 \addr_resp_reg[28]  ( .ip(n7522), .ck(clk), .q(N4216) );
  dp_1 \addr_resp_reg[29]  ( .ip(n7504), .ck(clk), .q(N4213) );
  dp_1 \addr_resp_reg[30]  ( .ip(n7486), .ck(clk), .q(N4210) );
  dp_1 \addr_resp_reg[31]  ( .ip(n7468), .ck(clk), .q(N4207) );
  dp_1 \iCache_data_wr_reg[0]  ( .ip(n7450), .ck(clk), .q(iCache_data_wr[0])
         );
  dp_1 \iCache_data_wr_reg[1]  ( .ip(n7449), .ck(clk), .q(iCache_data_wr[1])
         );
  dp_1 \iCache_data_wr_reg[2]  ( .ip(n7448), .ck(clk), .q(iCache_data_wr[2])
         );
  dp_1 \iCache_data_wr_reg[3]  ( .ip(n7447), .ck(clk), .q(iCache_data_wr[3])
         );
  dp_1 \iCache_data_wr_reg[4]  ( .ip(n7446), .ck(clk), .q(iCache_data_wr[4])
         );
  dp_1 \iCache_data_wr_reg[5]  ( .ip(n7445), .ck(clk), .q(iCache_data_wr[5])
         );
  dp_1 \iCache_data_wr_reg[6]  ( .ip(n7444), .ck(clk), .q(iCache_data_wr[6])
         );
  dp_1 \iCache_data_wr_reg[7]  ( .ip(n7443), .ck(clk), .q(iCache_data_wr[7])
         );
  dp_1 \iCache_data_wr_reg[8]  ( .ip(n7442), .ck(clk), .q(iCache_data_wr[8])
         );
  dp_1 \iCache_data_wr_reg[9]  ( .ip(n7441), .ck(clk), .q(iCache_data_wr[9])
         );
  dp_1 \iCache_data_wr_reg[10]  ( .ip(n7440), .ck(clk), .q(iCache_data_wr[10])
         );
  dp_1 \iCache_data_wr_reg[11]  ( .ip(n7439), .ck(clk), .q(iCache_data_wr[11])
         );
  dp_1 \iCache_data_wr_reg[12]  ( .ip(n7438), .ck(clk), .q(iCache_data_wr[12])
         );
  dp_1 \iCache_data_wr_reg[13]  ( .ip(n7437), .ck(clk), .q(iCache_data_wr[13])
         );
  dp_1 \iCache_data_wr_reg[14]  ( .ip(n7436), .ck(clk), .q(iCache_data_wr[14])
         );
  dp_1 \iCache_data_wr_reg[15]  ( .ip(n7435), .ck(clk), .q(iCache_data_wr[15])
         );
  dp_1 \iCache_data_wr_reg[16]  ( .ip(n7434), .ck(clk), .q(iCache_data_wr[16])
         );
  dp_1 \iCache_data_wr_reg[17]  ( .ip(n7433), .ck(clk), .q(iCache_data_wr[17])
         );
  dp_1 \iCache_data_wr_reg[18]  ( .ip(n7432), .ck(clk), .q(iCache_data_wr[18])
         );
  dp_1 \iCache_data_wr_reg[19]  ( .ip(n7431), .ck(clk), .q(iCache_data_wr[19])
         );
  dp_1 \iCache_data_wr_reg[20]  ( .ip(n7430), .ck(clk), .q(iCache_data_wr[20])
         );
  dp_1 \iCache_data_wr_reg[21]  ( .ip(n7429), .ck(clk), .q(iCache_data_wr[21])
         );
  dp_1 \iCache_data_wr_reg[22]  ( .ip(n7428), .ck(clk), .q(iCache_data_wr[22])
         );
  dp_1 \iCache_data_wr_reg[23]  ( .ip(n7427), .ck(clk), .q(iCache_data_wr[23])
         );
  dp_1 \iCache_data_wr_reg[24]  ( .ip(n7426), .ck(clk), .q(iCache_data_wr[24])
         );
  dp_1 \iCache_data_wr_reg[25]  ( .ip(n7425), .ck(clk), .q(iCache_data_wr[25])
         );
  dp_1 \iCache_data_wr_reg[26]  ( .ip(n7424), .ck(clk), .q(iCache_data_wr[26])
         );
  dp_1 \iCache_data_wr_reg[27]  ( .ip(n7423), .ck(clk), .q(iCache_data_wr[27])
         );
  dp_1 \iCache_data_wr_reg[28]  ( .ip(n7422), .ck(clk), .q(iCache_data_wr[28])
         );
  dp_1 \iCache_data_wr_reg[29]  ( .ip(n7421), .ck(clk), .q(iCache_data_wr[29])
         );
  dp_1 \iCache_data_wr_reg[30]  ( .ip(n7420), .ck(clk), .q(iCache_data_wr[30])
         );
  dp_1 \iCache_data_wr_reg[31]  ( .ip(n7419), .ck(clk), .q(iCache_data_wr[31])
         );
  dp_1 \cache_line_count_reg[0]  ( .ip(n7924), .ck(clk), .q(
        cache_line_count[0]) );
  dp_1 \cache_line_count_reg[1]  ( .ip(n7923), .ck(clk), .q(
        cache_line_count[1]) );
  dp_1 \cache_line_count_reg[2]  ( .ip(n7922), .ck(clk), .q(
        cache_line_count[2]) );
  dp_1 \cache_line_count_reg[3]  ( .ip(n7921), .ck(clk), .q(
        cache_line_count[3]) );
  dp_1 \cache_line_count_reg[4]  ( .ip(n7920), .ck(clk), .q(
        cache_line_count[4]) );
  dp_1 \cache_line_count_reg[5]  ( .ip(n7919), .ck(clk), .q(
        cache_line_count[5]) );
  dp_1 \cache_line_count_reg[6]  ( .ip(n7918), .ck(clk), .q(
        cache_line_count[6]) );
  dp_1 \cache_line_count_reg[7]  ( .ip(n7917), .ck(clk), .q(
        cache_line_count[7]) );
  dp_1 \cache_tag_B_reg[0][0]  ( .ip(n7890), .ck(clk), .q(\cache_tag_B[0][0] )
         );
  dp_1 \cache_tag_B_reg[0][1]  ( .ip(n7872), .ck(clk), .q(\cache_tag_B[0][1] )
         );
  dp_1 \cache_tag_B_reg[0][2]  ( .ip(n7854), .ck(clk), .q(\cache_tag_B[0][2] )
         );
  dp_1 \cache_tag_B_reg[0][3]  ( .ip(n7836), .ck(clk), .q(\cache_tag_B[0][3] )
         );
  dp_1 \cache_tag_B_reg[0][4]  ( .ip(n7818), .ck(clk), .q(\cache_tag_B[0][4] )
         );
  dp_1 \cache_tag_B_reg[0][5]  ( .ip(n7800), .ck(clk), .q(\cache_tag_B[0][5] )
         );
  dp_1 \cache_tag_B_reg[0][6]  ( .ip(n7782), .ck(clk), .q(\cache_tag_B[0][6] )
         );
  dp_1 \cache_tag_B_reg[0][7]  ( .ip(n7764), .ck(clk), .q(\cache_tag_B[0][7] )
         );
  dp_1 \cache_tag_B_reg[0][8]  ( .ip(n7746), .ck(clk), .q(\cache_tag_B[0][8] )
         );
  dp_1 \cache_tag_B_reg[0][9]  ( .ip(n7728), .ck(clk), .q(\cache_tag_B[0][9] )
         );
  dp_1 \cache_tag_B_reg[0][10]  ( .ip(n7710), .ck(clk), .q(
        \cache_tag_B[0][10] ) );
  dp_1 \cache_tag_B_reg[0][11]  ( .ip(n7692), .ck(clk), .q(
        \cache_tag_B[0][11] ) );
  dp_1 \cache_tag_B_reg[0][12]  ( .ip(n7674), .ck(clk), .q(
        \cache_tag_B[0][12] ) );
  dp_1 \cache_tag_B_reg[0][13]  ( .ip(n7656), .ck(clk), .q(
        \cache_tag_B[0][13] ) );
  dp_1 \cache_tag_B_reg[0][14]  ( .ip(n7638), .ck(clk), .q(
        \cache_tag_B[0][14] ) );
  dp_1 \cache_tag_B_reg[0][15]  ( .ip(n7620), .ck(clk), .q(
        \cache_tag_B[0][15] ) );
  dp_1 \cache_tag_B_reg[0][16]  ( .ip(n7602), .ck(clk), .q(
        \cache_tag_B[0][16] ) );
  dp_1 \cache_tag_B_reg[0][17]  ( .ip(n7584), .ck(clk), .q(
        \cache_tag_B[0][17] ) );
  dp_1 \cache_tag_B_reg[0][18]  ( .ip(n7566), .ck(clk), .q(
        \cache_tag_B[0][18] ) );
  dp_1 \cache_tag_B_reg[0][19]  ( .ip(n7548), .ck(clk), .q(
        \cache_tag_B[0][19] ) );
  dp_1 \cache_tag_B_reg[0][20]  ( .ip(n7530), .ck(clk), .q(
        \cache_tag_B[0][20] ) );
  dp_1 \cache_tag_B_reg[0][21]  ( .ip(n7512), .ck(clk), .q(
        \cache_tag_B[0][21] ) );
  dp_1 \cache_tag_B_reg[0][22]  ( .ip(n7494), .ck(clk), .q(
        \cache_tag_B[0][22] ) );
  dp_1 \cache_tag_B_reg[0][23]  ( .ip(n7476), .ck(clk), .q(
        \cache_tag_B[0][23] ) );
  dp_1 \cache_tag_B_reg[0][24]  ( .ip(n7458), .ck(clk), .q(
        \cache_tag_B[0][24] ) );
  dp_1 \cache_tag_B_reg[1][0]  ( .ip(n7889), .ck(clk), .q(\cache_tag_B[1][0] )
         );
  dp_1 \cache_tag_B_reg[1][1]  ( .ip(n7871), .ck(clk), .q(\cache_tag_B[1][1] )
         );
  dp_1 \cache_tag_B_reg[1][2]  ( .ip(n7853), .ck(clk), .q(\cache_tag_B[1][2] )
         );
  dp_1 \cache_tag_B_reg[1][3]  ( .ip(n7835), .ck(clk), .q(\cache_tag_B[1][3] )
         );
  dp_1 \cache_tag_B_reg[1][4]  ( .ip(n7817), .ck(clk), .q(\cache_tag_B[1][4] )
         );
  dp_1 \cache_tag_B_reg[1][5]  ( .ip(n7799), .ck(clk), .q(\cache_tag_B[1][5] )
         );
  dp_1 \cache_tag_B_reg[1][6]  ( .ip(n7781), .ck(clk), .q(\cache_tag_B[1][6] )
         );
  dp_1 \cache_tag_B_reg[1][7]  ( .ip(n7763), .ck(clk), .q(\cache_tag_B[1][7] )
         );
  dp_1 \cache_tag_B_reg[1][8]  ( .ip(n7745), .ck(clk), .q(\cache_tag_B[1][8] )
         );
  dp_1 \cache_tag_B_reg[1][9]  ( .ip(n7727), .ck(clk), .q(\cache_tag_B[1][9] )
         );
  dp_1 \cache_tag_B_reg[1][10]  ( .ip(n7709), .ck(clk), .q(
        \cache_tag_B[1][10] ) );
  dp_1 \cache_tag_B_reg[1][11]  ( .ip(n7691), .ck(clk), .q(
        \cache_tag_B[1][11] ) );
  dp_1 \cache_tag_B_reg[1][12]  ( .ip(n7673), .ck(clk), .q(
        \cache_tag_B[1][12] ) );
  dp_1 \cache_tag_B_reg[1][13]  ( .ip(n7655), .ck(clk), .q(
        \cache_tag_B[1][13] ) );
  dp_1 \cache_tag_B_reg[1][14]  ( .ip(n7637), .ck(clk), .q(
        \cache_tag_B[1][14] ) );
  dp_1 \cache_tag_B_reg[1][15]  ( .ip(n7619), .ck(clk), .q(
        \cache_tag_B[1][15] ) );
  dp_1 \cache_tag_B_reg[1][16]  ( .ip(n7601), .ck(clk), .q(
        \cache_tag_B[1][16] ) );
  dp_1 \cache_tag_B_reg[1][17]  ( .ip(n7583), .ck(clk), .q(
        \cache_tag_B[1][17] ) );
  dp_1 \cache_tag_B_reg[1][18]  ( .ip(n7565), .ck(clk), .q(
        \cache_tag_B[1][18] ) );
  dp_1 \cache_tag_B_reg[1][19]  ( .ip(n7547), .ck(clk), .q(
        \cache_tag_B[1][19] ) );
  dp_1 \cache_tag_B_reg[1][20]  ( .ip(n7529), .ck(clk), .q(
        \cache_tag_B[1][20] ) );
  dp_1 \cache_tag_B_reg[1][21]  ( .ip(n7511), .ck(clk), .q(
        \cache_tag_B[1][21] ) );
  dp_1 \cache_tag_B_reg[1][22]  ( .ip(n7493), .ck(clk), .q(
        \cache_tag_B[1][22] ) );
  dp_1 \cache_tag_B_reg[1][23]  ( .ip(n7475), .ck(clk), .q(
        \cache_tag_B[1][23] ) );
  dp_1 \cache_tag_B_reg[1][24]  ( .ip(n7457), .ck(clk), .q(
        \cache_tag_B[1][24] ) );
  dp_1 \cache_tag_B_reg[2][0]  ( .ip(n7888), .ck(clk), .q(\cache_tag_B[2][0] )
         );
  dp_1 \cache_tag_B_reg[2][1]  ( .ip(n7870), .ck(clk), .q(\cache_tag_B[2][1] )
         );
  dp_1 \cache_tag_B_reg[2][2]  ( .ip(n7852), .ck(clk), .q(\cache_tag_B[2][2] )
         );
  dp_1 \cache_tag_B_reg[2][3]  ( .ip(n7834), .ck(clk), .q(\cache_tag_B[2][3] )
         );
  dp_1 \cache_tag_B_reg[2][4]  ( .ip(n7816), .ck(clk), .q(\cache_tag_B[2][4] )
         );
  dp_1 \cache_tag_B_reg[2][5]  ( .ip(n7798), .ck(clk), .q(\cache_tag_B[2][5] )
         );
  dp_1 \cache_tag_B_reg[2][6]  ( .ip(n7780), .ck(clk), .q(\cache_tag_B[2][6] )
         );
  dp_1 \cache_tag_B_reg[2][7]  ( .ip(n7762), .ck(clk), .q(\cache_tag_B[2][7] )
         );
  dp_1 \cache_tag_B_reg[2][8]  ( .ip(n7744), .ck(clk), .q(\cache_tag_B[2][8] )
         );
  dp_1 \cache_tag_B_reg[2][9]  ( .ip(n7726), .ck(clk), .q(\cache_tag_B[2][9] )
         );
  dp_1 \cache_tag_B_reg[2][10]  ( .ip(n7708), .ck(clk), .q(
        \cache_tag_B[2][10] ) );
  dp_1 \cache_tag_B_reg[2][11]  ( .ip(n7690), .ck(clk), .q(
        \cache_tag_B[2][11] ) );
  dp_1 \cache_tag_B_reg[2][12]  ( .ip(n7672), .ck(clk), .q(
        \cache_tag_B[2][12] ) );
  dp_1 \cache_tag_B_reg[2][13]  ( .ip(n7654), .ck(clk), .q(
        \cache_tag_B[2][13] ) );
  dp_1 \cache_tag_B_reg[2][14]  ( .ip(n7636), .ck(clk), .q(
        \cache_tag_B[2][14] ) );
  dp_1 \cache_tag_B_reg[2][15]  ( .ip(n7618), .ck(clk), .q(
        \cache_tag_B[2][15] ) );
  dp_1 \cache_tag_B_reg[2][16]  ( .ip(n7600), .ck(clk), .q(
        \cache_tag_B[2][16] ) );
  dp_1 \cache_tag_B_reg[2][17]  ( .ip(n7582), .ck(clk), .q(
        \cache_tag_B[2][17] ) );
  dp_1 \cache_tag_B_reg[2][18]  ( .ip(n7564), .ck(clk), .q(
        \cache_tag_B[2][18] ) );
  dp_1 \cache_tag_B_reg[2][19]  ( .ip(n7546), .ck(clk), .q(
        \cache_tag_B[2][19] ) );
  dp_1 \cache_tag_B_reg[2][20]  ( .ip(n7528), .ck(clk), .q(
        \cache_tag_B[2][20] ) );
  dp_1 \cache_tag_B_reg[2][21]  ( .ip(n7510), .ck(clk), .q(
        \cache_tag_B[2][21] ) );
  dp_1 \cache_tag_B_reg[2][22]  ( .ip(n7492), .ck(clk), .q(
        \cache_tag_B[2][22] ) );
  dp_1 \cache_tag_B_reg[2][23]  ( .ip(n7474), .ck(clk), .q(
        \cache_tag_B[2][23] ) );
  dp_1 \cache_tag_B_reg[2][24]  ( .ip(n7456), .ck(clk), .q(
        \cache_tag_B[2][24] ) );
  dp_1 \cache_tag_B_reg[3][0]  ( .ip(n7887), .ck(clk), .q(\cache_tag_B[3][0] )
         );
  dp_1 \cache_tag_B_reg[3][1]  ( .ip(n7869), .ck(clk), .q(\cache_tag_B[3][1] )
         );
  dp_1 \cache_tag_B_reg[3][2]  ( .ip(n7851), .ck(clk), .q(\cache_tag_B[3][2] )
         );
  dp_1 \cache_tag_B_reg[3][3]  ( .ip(n7833), .ck(clk), .q(\cache_tag_B[3][3] )
         );
  dp_1 \cache_tag_B_reg[3][4]  ( .ip(n7815), .ck(clk), .q(\cache_tag_B[3][4] )
         );
  dp_1 \cache_tag_B_reg[3][5]  ( .ip(n7797), .ck(clk), .q(\cache_tag_B[3][5] )
         );
  dp_1 \cache_tag_B_reg[3][6]  ( .ip(n7779), .ck(clk), .q(\cache_tag_B[3][6] )
         );
  dp_1 \cache_tag_B_reg[3][7]  ( .ip(n7761), .ck(clk), .q(\cache_tag_B[3][7] )
         );
  dp_1 \cache_tag_B_reg[3][8]  ( .ip(n7743), .ck(clk), .q(\cache_tag_B[3][8] )
         );
  dp_1 \cache_tag_B_reg[3][9]  ( .ip(n7725), .ck(clk), .q(\cache_tag_B[3][9] )
         );
  dp_1 \cache_tag_B_reg[3][10]  ( .ip(n7707), .ck(clk), .q(
        \cache_tag_B[3][10] ) );
  dp_1 \cache_tag_B_reg[3][11]  ( .ip(n7689), .ck(clk), .q(
        \cache_tag_B[3][11] ) );
  dp_1 \cache_tag_B_reg[3][12]  ( .ip(n7671), .ck(clk), .q(
        \cache_tag_B[3][12] ) );
  dp_1 \cache_tag_B_reg[3][13]  ( .ip(n7653), .ck(clk), .q(
        \cache_tag_B[3][13] ) );
  dp_1 \cache_tag_B_reg[3][14]  ( .ip(n7635), .ck(clk), .q(
        \cache_tag_B[3][14] ) );
  dp_1 \cache_tag_B_reg[3][15]  ( .ip(n7617), .ck(clk), .q(
        \cache_tag_B[3][15] ) );
  dp_1 \cache_tag_B_reg[3][16]  ( .ip(n7599), .ck(clk), .q(
        \cache_tag_B[3][16] ) );
  dp_1 \cache_tag_B_reg[3][17]  ( .ip(n7581), .ck(clk), .q(
        \cache_tag_B[3][17] ) );
  dp_1 \cache_tag_B_reg[3][18]  ( .ip(n7563), .ck(clk), .q(
        \cache_tag_B[3][18] ) );
  dp_1 \cache_tag_B_reg[3][19]  ( .ip(n7545), .ck(clk), .q(
        \cache_tag_B[3][19] ) );
  dp_1 \cache_tag_B_reg[3][20]  ( .ip(n7527), .ck(clk), .q(
        \cache_tag_B[3][20] ) );
  dp_1 \cache_tag_B_reg[3][21]  ( .ip(n7509), .ck(clk), .q(
        \cache_tag_B[3][21] ) );
  dp_1 \cache_tag_B_reg[3][22]  ( .ip(n7491), .ck(clk), .q(
        \cache_tag_B[3][22] ) );
  dp_1 \cache_tag_B_reg[3][23]  ( .ip(n7473), .ck(clk), .q(
        \cache_tag_B[3][23] ) );
  dp_1 \cache_tag_B_reg[3][24]  ( .ip(n7455), .ck(clk), .q(
        \cache_tag_B[3][24] ) );
  dp_1 \cache_tag_B_reg[4][0]  ( .ip(n7886), .ck(clk), .q(\cache_tag_B[4][0] )
         );
  dp_1 \cache_tag_B_reg[4][1]  ( .ip(n7868), .ck(clk), .q(\cache_tag_B[4][1] )
         );
  dp_1 \cache_tag_B_reg[4][2]  ( .ip(n7850), .ck(clk), .q(\cache_tag_B[4][2] )
         );
  dp_1 \cache_tag_B_reg[4][3]  ( .ip(n7832), .ck(clk), .q(\cache_tag_B[4][3] )
         );
  dp_1 \cache_tag_B_reg[4][4]  ( .ip(n7814), .ck(clk), .q(\cache_tag_B[4][4] )
         );
  dp_1 \cache_tag_B_reg[4][5]  ( .ip(n7796), .ck(clk), .q(\cache_tag_B[4][5] )
         );
  dp_1 \cache_tag_B_reg[4][6]  ( .ip(n7778), .ck(clk), .q(\cache_tag_B[4][6] )
         );
  dp_1 \cache_tag_B_reg[4][7]  ( .ip(n7760), .ck(clk), .q(\cache_tag_B[4][7] )
         );
  dp_1 \cache_tag_B_reg[4][8]  ( .ip(n7742), .ck(clk), .q(\cache_tag_B[4][8] )
         );
  dp_1 \cache_tag_B_reg[4][9]  ( .ip(n7724), .ck(clk), .q(\cache_tag_B[4][9] )
         );
  dp_1 \cache_tag_B_reg[4][10]  ( .ip(n7706), .ck(clk), .q(
        \cache_tag_B[4][10] ) );
  dp_1 \cache_tag_B_reg[4][11]  ( .ip(n7688), .ck(clk), .q(
        \cache_tag_B[4][11] ) );
  dp_1 \cache_tag_B_reg[4][12]  ( .ip(n7670), .ck(clk), .q(
        \cache_tag_B[4][12] ) );
  dp_1 \cache_tag_B_reg[4][13]  ( .ip(n7652), .ck(clk), .q(
        \cache_tag_B[4][13] ) );
  dp_1 \cache_tag_B_reg[4][14]  ( .ip(n7634), .ck(clk), .q(
        \cache_tag_B[4][14] ) );
  dp_1 \cache_tag_B_reg[4][15]  ( .ip(n7616), .ck(clk), .q(
        \cache_tag_B[4][15] ) );
  dp_1 \cache_tag_B_reg[4][16]  ( .ip(n7598), .ck(clk), .q(
        \cache_tag_B[4][16] ) );
  dp_1 \cache_tag_B_reg[4][17]  ( .ip(n7580), .ck(clk), .q(
        \cache_tag_B[4][17] ) );
  dp_1 \cache_tag_B_reg[4][18]  ( .ip(n7562), .ck(clk), .q(
        \cache_tag_B[4][18] ) );
  dp_1 \cache_tag_B_reg[4][19]  ( .ip(n7544), .ck(clk), .q(
        \cache_tag_B[4][19] ) );
  dp_1 \cache_tag_B_reg[4][20]  ( .ip(n7526), .ck(clk), .q(
        \cache_tag_B[4][20] ) );
  dp_1 \cache_tag_B_reg[4][21]  ( .ip(n7508), .ck(clk), .q(
        \cache_tag_B[4][21] ) );
  dp_1 \cache_tag_B_reg[4][22]  ( .ip(n7490), .ck(clk), .q(
        \cache_tag_B[4][22] ) );
  dp_1 \cache_tag_B_reg[4][23]  ( .ip(n7472), .ck(clk), .q(
        \cache_tag_B[4][23] ) );
  dp_1 \cache_tag_B_reg[4][24]  ( .ip(n7454), .ck(clk), .q(
        \cache_tag_B[4][24] ) );
  dp_1 \cache_tag_B_reg[5][0]  ( .ip(n7885), .ck(clk), .q(\cache_tag_B[5][0] )
         );
  dp_1 \cache_tag_B_reg[5][1]  ( .ip(n7867), .ck(clk), .q(\cache_tag_B[5][1] )
         );
  dp_1 \cache_tag_B_reg[5][2]  ( .ip(n7849), .ck(clk), .q(\cache_tag_B[5][2] )
         );
  dp_1 \cache_tag_B_reg[5][3]  ( .ip(n7831), .ck(clk), .q(\cache_tag_B[5][3] )
         );
  dp_1 \cache_tag_B_reg[5][4]  ( .ip(n7813), .ck(clk), .q(\cache_tag_B[5][4] )
         );
  dp_1 \cache_tag_B_reg[5][5]  ( .ip(n7795), .ck(clk), .q(\cache_tag_B[5][5] )
         );
  dp_1 \cache_tag_B_reg[5][6]  ( .ip(n7777), .ck(clk), .q(\cache_tag_B[5][6] )
         );
  dp_1 \cache_tag_B_reg[5][7]  ( .ip(n7759), .ck(clk), .q(\cache_tag_B[5][7] )
         );
  dp_1 \cache_tag_B_reg[5][8]  ( .ip(n7741), .ck(clk), .q(\cache_tag_B[5][8] )
         );
  dp_1 \cache_tag_B_reg[5][9]  ( .ip(n7723), .ck(clk), .q(\cache_tag_B[5][9] )
         );
  dp_1 \cache_tag_B_reg[5][10]  ( .ip(n7705), .ck(clk), .q(
        \cache_tag_B[5][10] ) );
  dp_1 \cache_tag_B_reg[5][11]  ( .ip(n7687), .ck(clk), .q(
        \cache_tag_B[5][11] ) );
  dp_1 \cache_tag_B_reg[5][12]  ( .ip(n7669), .ck(clk), .q(
        \cache_tag_B[5][12] ) );
  dp_1 \cache_tag_B_reg[5][13]  ( .ip(n7651), .ck(clk), .q(
        \cache_tag_B[5][13] ) );
  dp_1 \cache_tag_B_reg[5][14]  ( .ip(n7633), .ck(clk), .q(
        \cache_tag_B[5][14] ) );
  dp_1 \cache_tag_B_reg[5][15]  ( .ip(n7615), .ck(clk), .q(
        \cache_tag_B[5][15] ) );
  dp_1 \cache_tag_B_reg[5][16]  ( .ip(n7597), .ck(clk), .q(
        \cache_tag_B[5][16] ) );
  dp_1 \cache_tag_B_reg[5][17]  ( .ip(n7579), .ck(clk), .q(
        \cache_tag_B[5][17] ) );
  dp_1 \cache_tag_B_reg[5][18]  ( .ip(n7561), .ck(clk), .q(
        \cache_tag_B[5][18] ) );
  dp_1 \cache_tag_B_reg[5][19]  ( .ip(n7543), .ck(clk), .q(
        \cache_tag_B[5][19] ) );
  dp_1 \cache_tag_B_reg[5][20]  ( .ip(n7525), .ck(clk), .q(
        \cache_tag_B[5][20] ) );
  dp_1 \cache_tag_B_reg[5][21]  ( .ip(n7507), .ck(clk), .q(
        \cache_tag_B[5][21] ) );
  dp_1 \cache_tag_B_reg[5][22]  ( .ip(n7489), .ck(clk), .q(
        \cache_tag_B[5][22] ) );
  dp_1 \cache_tag_B_reg[5][23]  ( .ip(n7471), .ck(clk), .q(
        \cache_tag_B[5][23] ) );
  dp_1 \cache_tag_B_reg[5][24]  ( .ip(n7453), .ck(clk), .q(
        \cache_tag_B[5][24] ) );
  dp_1 \cache_tag_B_reg[6][0]  ( .ip(n7884), .ck(clk), .q(\cache_tag_B[6][0] )
         );
  dp_1 \cache_tag_B_reg[6][1]  ( .ip(n7866), .ck(clk), .q(\cache_tag_B[6][1] )
         );
  dp_1 \cache_tag_B_reg[6][2]  ( .ip(n7848), .ck(clk), .q(\cache_tag_B[6][2] )
         );
  dp_1 \cache_tag_B_reg[6][3]  ( .ip(n7830), .ck(clk), .q(\cache_tag_B[6][3] )
         );
  dp_1 \cache_tag_B_reg[6][4]  ( .ip(n7812), .ck(clk), .q(\cache_tag_B[6][4] )
         );
  dp_1 \cache_tag_B_reg[6][5]  ( .ip(n7794), .ck(clk), .q(\cache_tag_B[6][5] )
         );
  dp_1 \cache_tag_B_reg[6][6]  ( .ip(n7776), .ck(clk), .q(\cache_tag_B[6][6] )
         );
  dp_1 \cache_tag_B_reg[6][7]  ( .ip(n7758), .ck(clk), .q(\cache_tag_B[6][7] )
         );
  dp_1 \cache_tag_B_reg[6][8]  ( .ip(n7740), .ck(clk), .q(\cache_tag_B[6][8] )
         );
  dp_1 \cache_tag_B_reg[6][9]  ( .ip(n7722), .ck(clk), .q(\cache_tag_B[6][9] )
         );
  dp_1 \cache_tag_B_reg[6][10]  ( .ip(n7704), .ck(clk), .q(
        \cache_tag_B[6][10] ) );
  dp_1 \cache_tag_B_reg[6][11]  ( .ip(n7686), .ck(clk), .q(
        \cache_tag_B[6][11] ) );
  dp_1 \cache_tag_B_reg[6][12]  ( .ip(n7668), .ck(clk), .q(
        \cache_tag_B[6][12] ) );
  dp_1 \cache_tag_B_reg[6][13]  ( .ip(n7650), .ck(clk), .q(
        \cache_tag_B[6][13] ) );
  dp_1 \cache_tag_B_reg[6][14]  ( .ip(n7632), .ck(clk), .q(
        \cache_tag_B[6][14] ) );
  dp_1 \cache_tag_B_reg[6][15]  ( .ip(n7614), .ck(clk), .q(
        \cache_tag_B[6][15] ) );
  dp_1 \cache_tag_B_reg[6][16]  ( .ip(n7596), .ck(clk), .q(
        \cache_tag_B[6][16] ) );
  dp_1 \cache_tag_B_reg[6][17]  ( .ip(n7578), .ck(clk), .q(
        \cache_tag_B[6][17] ) );
  dp_1 \cache_tag_B_reg[6][18]  ( .ip(n7560), .ck(clk), .q(
        \cache_tag_B[6][18] ) );
  dp_1 \cache_tag_B_reg[6][19]  ( .ip(n7542), .ck(clk), .q(
        \cache_tag_B[6][19] ) );
  dp_1 \cache_tag_B_reg[6][20]  ( .ip(n7524), .ck(clk), .q(
        \cache_tag_B[6][20] ) );
  dp_1 \cache_tag_B_reg[6][21]  ( .ip(n7506), .ck(clk), .q(
        \cache_tag_B[6][21] ) );
  dp_1 \cache_tag_B_reg[6][22]  ( .ip(n7488), .ck(clk), .q(
        \cache_tag_B[6][22] ) );
  dp_1 \cache_tag_B_reg[6][23]  ( .ip(n7470), .ck(clk), .q(
        \cache_tag_B[6][23] ) );
  dp_1 \cache_tag_B_reg[6][24]  ( .ip(n7452), .ck(clk), .q(
        \cache_tag_B[6][24] ) );
  dp_1 \cache_tag_B_reg[7][0]  ( .ip(n7883), .ck(clk), .q(\cache_tag_B[7][0] )
         );
  dp_1 \cache_tag_B_reg[7][1]  ( .ip(n7865), .ck(clk), .q(\cache_tag_B[7][1] )
         );
  dp_1 \cache_tag_B_reg[7][2]  ( .ip(n7847), .ck(clk), .q(\cache_tag_B[7][2] )
         );
  dp_1 \cache_tag_B_reg[7][3]  ( .ip(n7829), .ck(clk), .q(\cache_tag_B[7][3] )
         );
  dp_1 \cache_tag_B_reg[7][4]  ( .ip(n7811), .ck(clk), .q(\cache_tag_B[7][4] )
         );
  dp_1 \cache_tag_B_reg[7][5]  ( .ip(n7793), .ck(clk), .q(\cache_tag_B[7][5] )
         );
  dp_1 \cache_tag_B_reg[7][6]  ( .ip(n7775), .ck(clk), .q(\cache_tag_B[7][6] )
         );
  dp_1 \cache_tag_B_reg[7][7]  ( .ip(n7757), .ck(clk), .q(\cache_tag_B[7][7] )
         );
  dp_1 \cache_tag_B_reg[7][8]  ( .ip(n7739), .ck(clk), .q(\cache_tag_B[7][8] )
         );
  dp_1 \cache_tag_B_reg[7][9]  ( .ip(n7721), .ck(clk), .q(\cache_tag_B[7][9] )
         );
  dp_1 \cache_tag_B_reg[7][10]  ( .ip(n7703), .ck(clk), .q(
        \cache_tag_B[7][10] ) );
  dp_1 \cache_tag_B_reg[7][11]  ( .ip(n7685), .ck(clk), .q(
        \cache_tag_B[7][11] ) );
  dp_1 \cache_tag_B_reg[7][12]  ( .ip(n7667), .ck(clk), .q(
        \cache_tag_B[7][12] ) );
  dp_1 \cache_tag_B_reg[7][13]  ( .ip(n7649), .ck(clk), .q(
        \cache_tag_B[7][13] ) );
  dp_1 \cache_tag_B_reg[7][14]  ( .ip(n7631), .ck(clk), .q(
        \cache_tag_B[7][14] ) );
  dp_1 \cache_tag_B_reg[7][15]  ( .ip(n7613), .ck(clk), .q(
        \cache_tag_B[7][15] ) );
  dp_1 \cache_tag_B_reg[7][16]  ( .ip(n7595), .ck(clk), .q(
        \cache_tag_B[7][16] ) );
  dp_1 \cache_tag_B_reg[7][17]  ( .ip(n7577), .ck(clk), .q(
        \cache_tag_B[7][17] ) );
  dp_1 \cache_tag_B_reg[7][18]  ( .ip(n7559), .ck(clk), .q(
        \cache_tag_B[7][18] ) );
  dp_1 \cache_tag_B_reg[7][19]  ( .ip(n7541), .ck(clk), .q(
        \cache_tag_B[7][19] ) );
  dp_1 \cache_tag_B_reg[7][20]  ( .ip(n7523), .ck(clk), .q(
        \cache_tag_B[7][20] ) );
  dp_1 \cache_tag_B_reg[7][21]  ( .ip(n7505), .ck(clk), .q(
        \cache_tag_B[7][21] ) );
  dp_1 \cache_tag_B_reg[7][22]  ( .ip(n7487), .ck(clk), .q(
        \cache_tag_B[7][22] ) );
  dp_1 \cache_tag_B_reg[7][23]  ( .ip(n7469), .ck(clk), .q(
        \cache_tag_B[7][23] ) );
  dp_1 \cache_tag_B_reg[7][24]  ( .ip(n7451), .ck(clk), .q(
        \cache_tag_B[7][24] ) );
  dp_1 \cache_tag_A_reg[0][0]  ( .ip(n7898), .ck(clk), .q(\cache_tag_A[0][0] )
         );
  dp_1 \cache_tag_A_reg[0][1]  ( .ip(n7880), .ck(clk), .q(\cache_tag_A[0][1] )
         );
  dp_1 \cache_tag_A_reg[0][2]  ( .ip(n7862), .ck(clk), .q(\cache_tag_A[0][2] )
         );
  dp_1 \cache_tag_A_reg[0][3]  ( .ip(n7844), .ck(clk), .q(\cache_tag_A[0][3] )
         );
  dp_1 \cache_tag_A_reg[0][4]  ( .ip(n7826), .ck(clk), .q(\cache_tag_A[0][4] )
         );
  dp_1 \cache_tag_A_reg[0][5]  ( .ip(n7808), .ck(clk), .q(\cache_tag_A[0][5] )
         );
  dp_1 \cache_tag_A_reg[0][6]  ( .ip(n7790), .ck(clk), .q(\cache_tag_A[0][6] )
         );
  dp_1 \cache_tag_A_reg[0][7]  ( .ip(n7772), .ck(clk), .q(\cache_tag_A[0][7] )
         );
  dp_1 \cache_tag_A_reg[0][8]  ( .ip(n7754), .ck(clk), .q(\cache_tag_A[0][8] )
         );
  dp_1 \cache_tag_A_reg[0][9]  ( .ip(n7736), .ck(clk), .q(\cache_tag_A[0][9] )
         );
  dp_1 \cache_tag_A_reg[0][10]  ( .ip(n7718), .ck(clk), .q(
        \cache_tag_A[0][10] ) );
  dp_1 \cache_tag_A_reg[0][11]  ( .ip(n7700), .ck(clk), .q(
        \cache_tag_A[0][11] ) );
  dp_1 \cache_tag_A_reg[0][12]  ( .ip(n7682), .ck(clk), .q(
        \cache_tag_A[0][12] ) );
  dp_1 \cache_tag_A_reg[0][13]  ( .ip(n7664), .ck(clk), .q(
        \cache_tag_A[0][13] ) );
  dp_1 \cache_tag_A_reg[0][14]  ( .ip(n7646), .ck(clk), .q(
        \cache_tag_A[0][14] ) );
  dp_1 \cache_tag_A_reg[0][15]  ( .ip(n7628), .ck(clk), .q(
        \cache_tag_A[0][15] ) );
  dp_1 \cache_tag_A_reg[0][16]  ( .ip(n7610), .ck(clk), .q(
        \cache_tag_A[0][16] ) );
  dp_1 \cache_tag_A_reg[0][17]  ( .ip(n7592), .ck(clk), .q(
        \cache_tag_A[0][17] ) );
  dp_1 \cache_tag_A_reg[0][18]  ( .ip(n7574), .ck(clk), .q(
        \cache_tag_A[0][18] ) );
  dp_1 \cache_tag_A_reg[0][19]  ( .ip(n7556), .ck(clk), .q(
        \cache_tag_A[0][19] ) );
  dp_1 \cache_tag_A_reg[0][20]  ( .ip(n7538), .ck(clk), .q(
        \cache_tag_A[0][20] ) );
  dp_1 \cache_tag_A_reg[0][21]  ( .ip(n7520), .ck(clk), .q(
        \cache_tag_A[0][21] ) );
  dp_1 \cache_tag_A_reg[0][22]  ( .ip(n7502), .ck(clk), .q(
        \cache_tag_A[0][22] ) );
  dp_1 \cache_tag_A_reg[0][23]  ( .ip(n7484), .ck(clk), .q(
        \cache_tag_A[0][23] ) );
  dp_1 \cache_tag_A_reg[0][24]  ( .ip(n7466), .ck(clk), .q(
        \cache_tag_A[0][24] ) );
  dp_1 \cache_tag_A_reg[1][0]  ( .ip(n7897), .ck(clk), .q(\cache_tag_A[1][0] )
         );
  dp_1 \cache_tag_A_reg[1][1]  ( .ip(n7879), .ck(clk), .q(\cache_tag_A[1][1] )
         );
  dp_1 \cache_tag_A_reg[1][2]  ( .ip(n7861), .ck(clk), .q(\cache_tag_A[1][2] )
         );
  dp_1 \cache_tag_A_reg[1][3]  ( .ip(n7843), .ck(clk), .q(\cache_tag_A[1][3] )
         );
  dp_1 \cache_tag_A_reg[1][4]  ( .ip(n7825), .ck(clk), .q(\cache_tag_A[1][4] )
         );
  dp_1 \cache_tag_A_reg[1][5]  ( .ip(n7807), .ck(clk), .q(\cache_tag_A[1][5] )
         );
  dp_1 \cache_tag_A_reg[1][6]  ( .ip(n7789), .ck(clk), .q(\cache_tag_A[1][6] )
         );
  dp_1 \cache_tag_A_reg[1][7]  ( .ip(n7771), .ck(clk), .q(\cache_tag_A[1][7] )
         );
  dp_1 \cache_tag_A_reg[1][8]  ( .ip(n7753), .ck(clk), .q(\cache_tag_A[1][8] )
         );
  dp_1 \cache_tag_A_reg[1][9]  ( .ip(n7735), .ck(clk), .q(\cache_tag_A[1][9] )
         );
  dp_1 \cache_tag_A_reg[1][10]  ( .ip(n7717), .ck(clk), .q(
        \cache_tag_A[1][10] ) );
  dp_1 \cache_tag_A_reg[1][11]  ( .ip(n7699), .ck(clk), .q(
        \cache_tag_A[1][11] ) );
  dp_1 \cache_tag_A_reg[1][12]  ( .ip(n7681), .ck(clk), .q(
        \cache_tag_A[1][12] ) );
  dp_1 \cache_tag_A_reg[1][13]  ( .ip(n7663), .ck(clk), .q(
        \cache_tag_A[1][13] ) );
  dp_1 \cache_tag_A_reg[1][14]  ( .ip(n7645), .ck(clk), .q(
        \cache_tag_A[1][14] ) );
  dp_1 \cache_tag_A_reg[1][15]  ( .ip(n7627), .ck(clk), .q(
        \cache_tag_A[1][15] ) );
  dp_1 \cache_tag_A_reg[1][16]  ( .ip(n7609), .ck(clk), .q(
        \cache_tag_A[1][16] ) );
  dp_1 \cache_tag_A_reg[1][17]  ( .ip(n7591), .ck(clk), .q(
        \cache_tag_A[1][17] ) );
  dp_1 \cache_tag_A_reg[1][18]  ( .ip(n7573), .ck(clk), .q(
        \cache_tag_A[1][18] ) );
  dp_1 \cache_tag_A_reg[1][19]  ( .ip(n7555), .ck(clk), .q(
        \cache_tag_A[1][19] ) );
  dp_1 \cache_tag_A_reg[1][20]  ( .ip(n7537), .ck(clk), .q(
        \cache_tag_A[1][20] ) );
  dp_1 \cache_tag_A_reg[1][21]  ( .ip(n7519), .ck(clk), .q(
        \cache_tag_A[1][21] ) );
  dp_1 \cache_tag_A_reg[1][22]  ( .ip(n7501), .ck(clk), .q(
        \cache_tag_A[1][22] ) );
  dp_1 \cache_tag_A_reg[1][23]  ( .ip(n7483), .ck(clk), .q(
        \cache_tag_A[1][23] ) );
  dp_1 \cache_tag_A_reg[1][24]  ( .ip(n7465), .ck(clk), .q(
        \cache_tag_A[1][24] ) );
  dp_1 \cache_tag_A_reg[2][0]  ( .ip(n7896), .ck(clk), .q(\cache_tag_A[2][0] )
         );
  dp_1 \cache_tag_A_reg[2][1]  ( .ip(n7878), .ck(clk), .q(\cache_tag_A[2][1] )
         );
  dp_1 \cache_tag_A_reg[2][2]  ( .ip(n7860), .ck(clk), .q(\cache_tag_A[2][2] )
         );
  dp_1 \cache_tag_A_reg[2][3]  ( .ip(n7842), .ck(clk), .q(\cache_tag_A[2][3] )
         );
  dp_1 \cache_tag_A_reg[2][4]  ( .ip(n7824), .ck(clk), .q(\cache_tag_A[2][4] )
         );
  dp_1 \cache_tag_A_reg[2][5]  ( .ip(n7806), .ck(clk), .q(\cache_tag_A[2][5] )
         );
  dp_1 \cache_tag_A_reg[2][6]  ( .ip(n7788), .ck(clk), .q(\cache_tag_A[2][6] )
         );
  dp_1 \cache_tag_A_reg[2][7]  ( .ip(n7770), .ck(clk), .q(\cache_tag_A[2][7] )
         );
  dp_1 \cache_tag_A_reg[2][8]  ( .ip(n7752), .ck(clk), .q(\cache_tag_A[2][8] )
         );
  dp_1 \cache_tag_A_reg[2][9]  ( .ip(n7734), .ck(clk), .q(\cache_tag_A[2][9] )
         );
  dp_1 \cache_tag_A_reg[2][10]  ( .ip(n7716), .ck(clk), .q(
        \cache_tag_A[2][10] ) );
  dp_1 \cache_tag_A_reg[2][11]  ( .ip(n7698), .ck(clk), .q(
        \cache_tag_A[2][11] ) );
  dp_1 \cache_tag_A_reg[2][12]  ( .ip(n7680), .ck(clk), .q(
        \cache_tag_A[2][12] ) );
  dp_1 \cache_tag_A_reg[2][13]  ( .ip(n7662), .ck(clk), .q(
        \cache_tag_A[2][13] ) );
  dp_1 \cache_tag_A_reg[2][14]  ( .ip(n7644), .ck(clk), .q(
        \cache_tag_A[2][14] ) );
  dp_1 \cache_tag_A_reg[2][15]  ( .ip(n7626), .ck(clk), .q(
        \cache_tag_A[2][15] ) );
  dp_1 \cache_tag_A_reg[2][16]  ( .ip(n7608), .ck(clk), .q(
        \cache_tag_A[2][16] ) );
  dp_1 \cache_tag_A_reg[2][17]  ( .ip(n7590), .ck(clk), .q(
        \cache_tag_A[2][17] ) );
  dp_1 \cache_tag_A_reg[2][18]  ( .ip(n7572), .ck(clk), .q(
        \cache_tag_A[2][18] ) );
  dp_1 \cache_tag_A_reg[2][19]  ( .ip(n7554), .ck(clk), .q(
        \cache_tag_A[2][19] ) );
  dp_1 \cache_tag_A_reg[2][20]  ( .ip(n7536), .ck(clk), .q(
        \cache_tag_A[2][20] ) );
  dp_1 \cache_tag_A_reg[2][21]  ( .ip(n7518), .ck(clk), .q(
        \cache_tag_A[2][21] ) );
  dp_1 \cache_tag_A_reg[2][22]  ( .ip(n7500), .ck(clk), .q(
        \cache_tag_A[2][22] ) );
  dp_1 \cache_tag_A_reg[2][23]  ( .ip(n7482), .ck(clk), .q(
        \cache_tag_A[2][23] ) );
  dp_1 \cache_tag_A_reg[2][24]  ( .ip(n7464), .ck(clk), .q(
        \cache_tag_A[2][24] ) );
  dp_1 \cache_tag_A_reg[3][0]  ( .ip(n7895), .ck(clk), .q(\cache_tag_A[3][0] )
         );
  dp_1 \cache_tag_A_reg[3][1]  ( .ip(n7877), .ck(clk), .q(\cache_tag_A[3][1] )
         );
  dp_1 \cache_tag_A_reg[3][2]  ( .ip(n7859), .ck(clk), .q(\cache_tag_A[3][2] )
         );
  dp_1 \cache_tag_A_reg[3][3]  ( .ip(n7841), .ck(clk), .q(\cache_tag_A[3][3] )
         );
  dp_1 \cache_tag_A_reg[3][4]  ( .ip(n7823), .ck(clk), .q(\cache_tag_A[3][4] )
         );
  dp_1 \cache_tag_A_reg[3][5]  ( .ip(n7805), .ck(clk), .q(\cache_tag_A[3][5] )
         );
  dp_1 \cache_tag_A_reg[3][6]  ( .ip(n7787), .ck(clk), .q(\cache_tag_A[3][6] )
         );
  dp_1 \cache_tag_A_reg[3][7]  ( .ip(n7769), .ck(clk), .q(\cache_tag_A[3][7] )
         );
  dp_1 \cache_tag_A_reg[3][8]  ( .ip(n7751), .ck(clk), .q(\cache_tag_A[3][8] )
         );
  dp_1 \cache_tag_A_reg[3][9]  ( .ip(n7733), .ck(clk), .q(\cache_tag_A[3][9] )
         );
  dp_1 \cache_tag_A_reg[3][10]  ( .ip(n7715), .ck(clk), .q(
        \cache_tag_A[3][10] ) );
  dp_1 \cache_tag_A_reg[3][11]  ( .ip(n7697), .ck(clk), .q(
        \cache_tag_A[3][11] ) );
  dp_1 \cache_tag_A_reg[3][12]  ( .ip(n7679), .ck(clk), .q(
        \cache_tag_A[3][12] ) );
  dp_1 \cache_tag_A_reg[3][13]  ( .ip(n7661), .ck(clk), .q(
        \cache_tag_A[3][13] ) );
  dp_1 \cache_tag_A_reg[3][14]  ( .ip(n7643), .ck(clk), .q(
        \cache_tag_A[3][14] ) );
  dp_1 \cache_tag_A_reg[3][15]  ( .ip(n7625), .ck(clk), .q(
        \cache_tag_A[3][15] ) );
  dp_1 \cache_tag_A_reg[3][16]  ( .ip(n7607), .ck(clk), .q(
        \cache_tag_A[3][16] ) );
  dp_1 \cache_tag_A_reg[3][17]  ( .ip(n7589), .ck(clk), .q(
        \cache_tag_A[3][17] ) );
  dp_1 \cache_tag_A_reg[3][18]  ( .ip(n7571), .ck(clk), .q(
        \cache_tag_A[3][18] ) );
  dp_1 \cache_tag_A_reg[3][19]  ( .ip(n7553), .ck(clk), .q(
        \cache_tag_A[3][19] ) );
  dp_1 \cache_tag_A_reg[3][20]  ( .ip(n7535), .ck(clk), .q(
        \cache_tag_A[3][20] ) );
  dp_1 \cache_tag_A_reg[3][21]  ( .ip(n7517), .ck(clk), .q(
        \cache_tag_A[3][21] ) );
  dp_1 \cache_tag_A_reg[3][22]  ( .ip(n7499), .ck(clk), .q(
        \cache_tag_A[3][22] ) );
  dp_1 \cache_tag_A_reg[3][23]  ( .ip(n7481), .ck(clk), .q(
        \cache_tag_A[3][23] ) );
  dp_1 \cache_tag_A_reg[3][24]  ( .ip(n7463), .ck(clk), .q(
        \cache_tag_A[3][24] ) );
  dp_1 \cache_tag_A_reg[4][0]  ( .ip(n7894), .ck(clk), .q(\cache_tag_A[4][0] )
         );
  dp_1 \cache_tag_A_reg[4][1]  ( .ip(n7876), .ck(clk), .q(\cache_tag_A[4][1] )
         );
  dp_1 \cache_tag_A_reg[4][2]  ( .ip(n7858), .ck(clk), .q(\cache_tag_A[4][2] )
         );
  dp_1 \cache_tag_A_reg[4][3]  ( .ip(n7840), .ck(clk), .q(\cache_tag_A[4][3] )
         );
  dp_1 \cache_tag_A_reg[4][4]  ( .ip(n7822), .ck(clk), .q(\cache_tag_A[4][4] )
         );
  dp_1 \cache_tag_A_reg[4][5]  ( .ip(n7804), .ck(clk), .q(\cache_tag_A[4][5] )
         );
  dp_1 \cache_tag_A_reg[4][6]  ( .ip(n7786), .ck(clk), .q(\cache_tag_A[4][6] )
         );
  dp_1 \cache_tag_A_reg[4][7]  ( .ip(n7768), .ck(clk), .q(\cache_tag_A[4][7] )
         );
  dp_1 \cache_tag_A_reg[4][8]  ( .ip(n7750), .ck(clk), .q(\cache_tag_A[4][8] )
         );
  dp_1 \cache_tag_A_reg[4][9]  ( .ip(n7732), .ck(clk), .q(\cache_tag_A[4][9] )
         );
  dp_1 \cache_tag_A_reg[4][10]  ( .ip(n7714), .ck(clk), .q(
        \cache_tag_A[4][10] ) );
  dp_1 \cache_tag_A_reg[4][11]  ( .ip(n7696), .ck(clk), .q(
        \cache_tag_A[4][11] ) );
  dp_1 \cache_tag_A_reg[4][12]  ( .ip(n7678), .ck(clk), .q(
        \cache_tag_A[4][12] ) );
  dp_1 \cache_tag_A_reg[4][13]  ( .ip(n7660), .ck(clk), .q(
        \cache_tag_A[4][13] ) );
  dp_1 \cache_tag_A_reg[4][14]  ( .ip(n7642), .ck(clk), .q(
        \cache_tag_A[4][14] ) );
  dp_1 \cache_tag_A_reg[4][15]  ( .ip(n7624), .ck(clk), .q(
        \cache_tag_A[4][15] ) );
  dp_1 \cache_tag_A_reg[4][16]  ( .ip(n7606), .ck(clk), .q(
        \cache_tag_A[4][16] ) );
  dp_1 \cache_tag_A_reg[4][17]  ( .ip(n7588), .ck(clk), .q(
        \cache_tag_A[4][17] ) );
  dp_1 \cache_tag_A_reg[4][18]  ( .ip(n7570), .ck(clk), .q(
        \cache_tag_A[4][18] ) );
  dp_1 \cache_tag_A_reg[4][19]  ( .ip(n7552), .ck(clk), .q(
        \cache_tag_A[4][19] ) );
  dp_1 \cache_tag_A_reg[4][20]  ( .ip(n7534), .ck(clk), .q(
        \cache_tag_A[4][20] ) );
  dp_1 \cache_tag_A_reg[4][21]  ( .ip(n7516), .ck(clk), .q(
        \cache_tag_A[4][21] ) );
  dp_1 \cache_tag_A_reg[4][22]  ( .ip(n7498), .ck(clk), .q(
        \cache_tag_A[4][22] ) );
  dp_1 \cache_tag_A_reg[4][23]  ( .ip(n7480), .ck(clk), .q(
        \cache_tag_A[4][23] ) );
  dp_1 \cache_tag_A_reg[4][24]  ( .ip(n7462), .ck(clk), .q(
        \cache_tag_A[4][24] ) );
  dp_1 \cache_tag_A_reg[5][0]  ( .ip(n7893), .ck(clk), .q(\cache_tag_A[5][0] )
         );
  dp_1 \cache_tag_A_reg[5][1]  ( .ip(n7875), .ck(clk), .q(\cache_tag_A[5][1] )
         );
  dp_1 \cache_tag_A_reg[5][2]  ( .ip(n7857), .ck(clk), .q(\cache_tag_A[5][2] )
         );
  dp_1 \cache_tag_A_reg[5][3]  ( .ip(n7839), .ck(clk), .q(\cache_tag_A[5][3] )
         );
  dp_1 \cache_tag_A_reg[5][4]  ( .ip(n7821), .ck(clk), .q(\cache_tag_A[5][4] )
         );
  dp_1 \cache_tag_A_reg[5][5]  ( .ip(n7803), .ck(clk), .q(\cache_tag_A[5][5] )
         );
  dp_1 \cache_tag_A_reg[5][6]  ( .ip(n7785), .ck(clk), .q(\cache_tag_A[5][6] )
         );
  dp_1 \cache_tag_A_reg[5][7]  ( .ip(n7767), .ck(clk), .q(\cache_tag_A[5][7] )
         );
  dp_1 \cache_tag_A_reg[5][8]  ( .ip(n7749), .ck(clk), .q(\cache_tag_A[5][8] )
         );
  dp_1 \cache_tag_A_reg[5][9]  ( .ip(n7731), .ck(clk), .q(\cache_tag_A[5][9] )
         );
  dp_1 \cache_tag_A_reg[5][10]  ( .ip(n7713), .ck(clk), .q(
        \cache_tag_A[5][10] ) );
  dp_1 \cache_tag_A_reg[5][11]  ( .ip(n7695), .ck(clk), .q(
        \cache_tag_A[5][11] ) );
  dp_1 \cache_tag_A_reg[5][12]  ( .ip(n7677), .ck(clk), .q(
        \cache_tag_A[5][12] ) );
  dp_1 \cache_tag_A_reg[5][13]  ( .ip(n7659), .ck(clk), .q(
        \cache_tag_A[5][13] ) );
  dp_1 \cache_tag_A_reg[5][14]  ( .ip(n7641), .ck(clk), .q(
        \cache_tag_A[5][14] ) );
  dp_1 \cache_tag_A_reg[5][15]  ( .ip(n7623), .ck(clk), .q(
        \cache_tag_A[5][15] ) );
  dp_1 \cache_tag_A_reg[5][16]  ( .ip(n7605), .ck(clk), .q(
        \cache_tag_A[5][16] ) );
  dp_1 \cache_tag_A_reg[5][17]  ( .ip(n7587), .ck(clk), .q(
        \cache_tag_A[5][17] ) );
  dp_1 \cache_tag_A_reg[5][18]  ( .ip(n7569), .ck(clk), .q(
        \cache_tag_A[5][18] ) );
  dp_1 \cache_tag_A_reg[5][19]  ( .ip(n7551), .ck(clk), .q(
        \cache_tag_A[5][19] ) );
  dp_1 \cache_tag_A_reg[5][20]  ( .ip(n7533), .ck(clk), .q(
        \cache_tag_A[5][20] ) );
  dp_1 \cache_tag_A_reg[5][21]  ( .ip(n7515), .ck(clk), .q(
        \cache_tag_A[5][21] ) );
  dp_1 \cache_tag_A_reg[5][22]  ( .ip(n7497), .ck(clk), .q(
        \cache_tag_A[5][22] ) );
  dp_1 \cache_tag_A_reg[5][23]  ( .ip(n7479), .ck(clk), .q(
        \cache_tag_A[5][23] ) );
  dp_1 \cache_tag_A_reg[5][24]  ( .ip(n7461), .ck(clk), .q(
        \cache_tag_A[5][24] ) );
  dp_1 \cache_tag_A_reg[6][0]  ( .ip(n7892), .ck(clk), .q(\cache_tag_A[6][0] )
         );
  dp_1 \cache_tag_A_reg[6][1]  ( .ip(n7874), .ck(clk), .q(\cache_tag_A[6][1] )
         );
  dp_1 \cache_tag_A_reg[6][2]  ( .ip(n7856), .ck(clk), .q(\cache_tag_A[6][2] )
         );
  dp_1 \cache_tag_A_reg[6][3]  ( .ip(n7838), .ck(clk), .q(\cache_tag_A[6][3] )
         );
  dp_1 \cache_tag_A_reg[6][4]  ( .ip(n7820), .ck(clk), .q(\cache_tag_A[6][4] )
         );
  dp_1 \cache_tag_A_reg[6][5]  ( .ip(n7802), .ck(clk), .q(\cache_tag_A[6][5] )
         );
  dp_1 \cache_tag_A_reg[6][6]  ( .ip(n7784), .ck(clk), .q(\cache_tag_A[6][6] )
         );
  dp_1 \cache_tag_A_reg[6][7]  ( .ip(n7766), .ck(clk), .q(\cache_tag_A[6][7] )
         );
  dp_1 \cache_tag_A_reg[6][8]  ( .ip(n7748), .ck(clk), .q(\cache_tag_A[6][8] )
         );
  dp_1 \cache_tag_A_reg[6][9]  ( .ip(n7730), .ck(clk), .q(\cache_tag_A[6][9] )
         );
  dp_1 \cache_tag_A_reg[6][10]  ( .ip(n7712), .ck(clk), .q(
        \cache_tag_A[6][10] ) );
  dp_1 \cache_tag_A_reg[6][11]  ( .ip(n7694), .ck(clk), .q(
        \cache_tag_A[6][11] ) );
  dp_1 \cache_tag_A_reg[6][12]  ( .ip(n7676), .ck(clk), .q(
        \cache_tag_A[6][12] ) );
  dp_1 \cache_tag_A_reg[6][13]  ( .ip(n7658), .ck(clk), .q(
        \cache_tag_A[6][13] ) );
  dp_1 \cache_tag_A_reg[6][14]  ( .ip(n7640), .ck(clk), .q(
        \cache_tag_A[6][14] ) );
  dp_1 \cache_tag_A_reg[6][15]  ( .ip(n7622), .ck(clk), .q(
        \cache_tag_A[6][15] ) );
  dp_1 \cache_tag_A_reg[6][16]  ( .ip(n7604), .ck(clk), .q(
        \cache_tag_A[6][16] ) );
  dp_1 \cache_tag_A_reg[6][17]  ( .ip(n7586), .ck(clk), .q(
        \cache_tag_A[6][17] ) );
  dp_1 \cache_tag_A_reg[6][18]  ( .ip(n7568), .ck(clk), .q(
        \cache_tag_A[6][18] ) );
  dp_1 \cache_tag_A_reg[6][19]  ( .ip(n7550), .ck(clk), .q(
        \cache_tag_A[6][19] ) );
  dp_1 \cache_tag_A_reg[6][20]  ( .ip(n7532), .ck(clk), .q(
        \cache_tag_A[6][20] ) );
  dp_1 \cache_tag_A_reg[6][21]  ( .ip(n7514), .ck(clk), .q(
        \cache_tag_A[6][21] ) );
  dp_1 \cache_tag_A_reg[6][22]  ( .ip(n7496), .ck(clk), .q(
        \cache_tag_A[6][22] ) );
  dp_1 \cache_tag_A_reg[6][23]  ( .ip(n7478), .ck(clk), .q(
        \cache_tag_A[6][23] ) );
  dp_1 \cache_tag_A_reg[6][24]  ( .ip(n7460), .ck(clk), .q(
        \cache_tag_A[6][24] ) );
  dp_1 \cache_tag_A_reg[7][0]  ( .ip(n7891), .ck(clk), .q(\cache_tag_A[7][0] )
         );
  dp_1 \cache_tag_A_reg[7][1]  ( .ip(n7873), .ck(clk), .q(\cache_tag_A[7][1] )
         );
  dp_1 \cache_tag_A_reg[7][2]  ( .ip(n7855), .ck(clk), .q(\cache_tag_A[7][2] )
         );
  dp_1 \cache_tag_A_reg[7][3]  ( .ip(n7837), .ck(clk), .q(\cache_tag_A[7][3] )
         );
  dp_1 \cache_tag_A_reg[7][4]  ( .ip(n7819), .ck(clk), .q(\cache_tag_A[7][4] )
         );
  dp_1 \cache_tag_A_reg[7][5]  ( .ip(n7801), .ck(clk), .q(\cache_tag_A[7][5] )
         );
  dp_1 \cache_tag_A_reg[7][6]  ( .ip(n7783), .ck(clk), .q(\cache_tag_A[7][6] )
         );
  dp_1 \cache_tag_A_reg[7][7]  ( .ip(n7765), .ck(clk), .q(\cache_tag_A[7][7] )
         );
  dp_1 \cache_tag_A_reg[7][8]  ( .ip(n7747), .ck(clk), .q(\cache_tag_A[7][8] )
         );
  dp_1 \cache_tag_A_reg[7][9]  ( .ip(n7729), .ck(clk), .q(\cache_tag_A[7][9] )
         );
  dp_1 \cache_tag_A_reg[7][10]  ( .ip(n7711), .ck(clk), .q(
        \cache_tag_A[7][10] ) );
  dp_1 \cache_tag_A_reg[7][11]  ( .ip(n7693), .ck(clk), .q(
        \cache_tag_A[7][11] ) );
  dp_1 \cache_tag_A_reg[7][12]  ( .ip(n7675), .ck(clk), .q(
        \cache_tag_A[7][12] ) );
  dp_1 \cache_tag_A_reg[7][13]  ( .ip(n7657), .ck(clk), .q(
        \cache_tag_A[7][13] ) );
  dp_1 \cache_tag_A_reg[7][14]  ( .ip(n7639), .ck(clk), .q(
        \cache_tag_A[7][14] ) );
  dp_1 \cache_tag_A_reg[7][15]  ( .ip(n7621), .ck(clk), .q(
        \cache_tag_A[7][15] ) );
  dp_1 \cache_tag_A_reg[7][16]  ( .ip(n7603), .ck(clk), .q(
        \cache_tag_A[7][16] ) );
  dp_1 \cache_tag_A_reg[7][17]  ( .ip(n7585), .ck(clk), .q(
        \cache_tag_A[7][17] ) );
  dp_1 \cache_tag_A_reg[7][18]  ( .ip(n7567), .ck(clk), .q(
        \cache_tag_A[7][18] ) );
  dp_1 \cache_tag_A_reg[7][19]  ( .ip(n7549), .ck(clk), .q(
        \cache_tag_A[7][19] ) );
  dp_1 \cache_tag_A_reg[7][20]  ( .ip(n7531), .ck(clk), .q(
        \cache_tag_A[7][20] ) );
  dp_1 \cache_tag_A_reg[7][21]  ( .ip(n7513), .ck(clk), .q(
        \cache_tag_A[7][21] ) );
  dp_1 \cache_tag_A_reg[7][22]  ( .ip(n7495), .ck(clk), .q(
        \cache_tag_A[7][22] ) );
  dp_1 \cache_tag_A_reg[7][23]  ( .ip(n7477), .ck(clk), .q(
        \cache_tag_A[7][23] ) );
  dp_1 \cache_tag_A_reg[7][24]  ( .ip(n7459), .ck(clk), .q(
        \cache_tag_A[7][24] ) );
  dp_1 \cache_data_B_reg[0][0]  ( .ip(n6360), .ck(clk), .q(
        \cache_data_B[0][0] ) );
  dp_1 \cache_data_B_reg[0][1]  ( .ip(n6359), .ck(clk), .q(
        \cache_data_B[0][1] ) );
  dp_1 \cache_data_B_reg[0][2]  ( .ip(n6358), .ck(clk), .q(
        \cache_data_B[0][2] ) );
  dp_1 \cache_data_B_reg[0][3]  ( .ip(n6357), .ck(clk), .q(
        \cache_data_B[0][3] ) );
  dp_1 \cache_data_B_reg[0][4]  ( .ip(n6356), .ck(clk), .q(
        \cache_data_B[0][4] ) );
  dp_1 \cache_data_B_reg[0][5]  ( .ip(n6355), .ck(clk), .q(
        \cache_data_B[0][5] ) );
  dp_1 \cache_data_B_reg[0][6]  ( .ip(n6354), .ck(clk), .q(
        \cache_data_B[0][6] ) );
  dp_1 \cache_data_B_reg[0][7]  ( .ip(n6353), .ck(clk), .q(
        \cache_data_B[0][7] ) );
  dp_1 \cache_data_B_reg[0][8]  ( .ip(n6352), .ck(clk), .q(
        \cache_data_B[0][8] ) );
  dp_1 \cache_data_B_reg[0][9]  ( .ip(n6351), .ck(clk), .q(
        \cache_data_B[0][9] ) );
  dp_1 \cache_data_B_reg[0][10]  ( .ip(n6350), .ck(clk), .q(
        \cache_data_B[0][10] ) );
  dp_1 \cache_data_B_reg[0][11]  ( .ip(n6349), .ck(clk), .q(
        \cache_data_B[0][11] ) );
  dp_1 \cache_data_B_reg[0][12]  ( .ip(n6348), .ck(clk), .q(
        \cache_data_B[0][12] ) );
  dp_1 \cache_data_B_reg[0][13]  ( .ip(n6347), .ck(clk), .q(
        \cache_data_B[0][13] ) );
  dp_1 \cache_data_B_reg[0][14]  ( .ip(n6346), .ck(clk), .q(
        \cache_data_B[0][14] ) );
  dp_1 \cache_data_B_reg[0][15]  ( .ip(n6345), .ck(clk), .q(
        \cache_data_B[0][15] ) );
  dp_1 \cache_data_B_reg[0][16]  ( .ip(n6344), .ck(clk), .q(
        \cache_data_B[0][16] ) );
  dp_1 \cache_data_B_reg[0][17]  ( .ip(n6343), .ck(clk), .q(
        \cache_data_B[0][17] ) );
  dp_1 \cache_data_B_reg[0][18]  ( .ip(n6342), .ck(clk), .q(
        \cache_data_B[0][18] ) );
  dp_1 \cache_data_B_reg[0][19]  ( .ip(n6341), .ck(clk), .q(
        \cache_data_B[0][19] ) );
  dp_1 \cache_data_B_reg[0][20]  ( .ip(n6340), .ck(clk), .q(
        \cache_data_B[0][20] ) );
  dp_1 \cache_data_B_reg[0][21]  ( .ip(n6339), .ck(clk), .q(
        \cache_data_B[0][21] ) );
  dp_1 \cache_data_B_reg[0][22]  ( .ip(n6338), .ck(clk), .q(
        \cache_data_B[0][22] ) );
  dp_1 \cache_data_B_reg[0][23]  ( .ip(n6337), .ck(clk), .q(
        \cache_data_B[0][23] ) );
  dp_1 \cache_data_B_reg[0][24]  ( .ip(n6336), .ck(clk), .q(
        \cache_data_B[0][24] ) );
  dp_1 \cache_data_B_reg[0][25]  ( .ip(n6335), .ck(clk), .q(
        \cache_data_B[0][25] ) );
  dp_1 \cache_data_B_reg[0][26]  ( .ip(n6334), .ck(clk), .q(
        \cache_data_B[0][26] ) );
  dp_1 \cache_data_B_reg[0][27]  ( .ip(n6333), .ck(clk), .q(
        \cache_data_B[0][27] ) );
  dp_1 \cache_data_B_reg[0][28]  ( .ip(n6332), .ck(clk), .q(
        \cache_data_B[0][28] ) );
  dp_1 \cache_data_B_reg[0][29]  ( .ip(n6331), .ck(clk), .q(
        \cache_data_B[0][29] ) );
  dp_1 \cache_data_B_reg[0][30]  ( .ip(n6330), .ck(clk), .q(
        \cache_data_B[0][30] ) );
  dp_1 \cache_data_B_reg[0][31]  ( .ip(n6329), .ck(clk), .q(
        \cache_data_B[0][31] ) );
  dp_1 \cache_data_B_reg[1][0]  ( .ip(n6232), .ck(clk), .q(
        \cache_data_B[1][0] ) );
  dp_1 \cache_data_B_reg[1][1]  ( .ip(n6231), .ck(clk), .q(
        \cache_data_B[1][1] ) );
  dp_1 \cache_data_B_reg[1][2]  ( .ip(n6230), .ck(clk), .q(
        \cache_data_B[1][2] ) );
  dp_1 \cache_data_B_reg[1][3]  ( .ip(n6229), .ck(clk), .q(
        \cache_data_B[1][3] ) );
  dp_1 \cache_data_B_reg[1][4]  ( .ip(n6228), .ck(clk), .q(
        \cache_data_B[1][4] ) );
  dp_1 \cache_data_B_reg[1][5]  ( .ip(n6227), .ck(clk), .q(
        \cache_data_B[1][5] ) );
  dp_1 \cache_data_B_reg[1][6]  ( .ip(n6226), .ck(clk), .q(
        \cache_data_B[1][6] ) );
  dp_1 \cache_data_B_reg[1][7]  ( .ip(n6225), .ck(clk), .q(
        \cache_data_B[1][7] ) );
  dp_1 \cache_data_B_reg[1][8]  ( .ip(n6224), .ck(clk), .q(
        \cache_data_B[1][8] ) );
  dp_1 \cache_data_B_reg[1][9]  ( .ip(n6223), .ck(clk), .q(
        \cache_data_B[1][9] ) );
  dp_1 \cache_data_B_reg[1][10]  ( .ip(n6222), .ck(clk), .q(
        \cache_data_B[1][10] ) );
  dp_1 \cache_data_B_reg[1][11]  ( .ip(n6221), .ck(clk), .q(
        \cache_data_B[1][11] ) );
  dp_1 \cache_data_B_reg[1][12]  ( .ip(n6220), .ck(clk), .q(
        \cache_data_B[1][12] ) );
  dp_1 \cache_data_B_reg[1][13]  ( .ip(n6219), .ck(clk), .q(
        \cache_data_B[1][13] ) );
  dp_1 \cache_data_B_reg[1][14]  ( .ip(n6218), .ck(clk), .q(
        \cache_data_B[1][14] ) );
  dp_1 \cache_data_B_reg[1][15]  ( .ip(n6217), .ck(clk), .q(
        \cache_data_B[1][15] ) );
  dp_1 \cache_data_B_reg[1][16]  ( .ip(n6216), .ck(clk), .q(
        \cache_data_B[1][16] ) );
  dp_1 \cache_data_B_reg[1][17]  ( .ip(n6215), .ck(clk), .q(
        \cache_data_B[1][17] ) );
  dp_1 \cache_data_B_reg[1][18]  ( .ip(n6214), .ck(clk), .q(
        \cache_data_B[1][18] ) );
  dp_1 \cache_data_B_reg[1][19]  ( .ip(n6213), .ck(clk), .q(
        \cache_data_B[1][19] ) );
  dp_1 \cache_data_B_reg[1][20]  ( .ip(n6212), .ck(clk), .q(
        \cache_data_B[1][20] ) );
  dp_1 \cache_data_B_reg[1][21]  ( .ip(n6211), .ck(clk), .q(
        \cache_data_B[1][21] ) );
  dp_1 \cache_data_B_reg[1][22]  ( .ip(n6210), .ck(clk), .q(
        \cache_data_B[1][22] ) );
  dp_1 \cache_data_B_reg[1][23]  ( .ip(n6209), .ck(clk), .q(
        \cache_data_B[1][23] ) );
  dp_1 \cache_data_B_reg[1][24]  ( .ip(n6208), .ck(clk), .q(
        \cache_data_B[1][24] ) );
  dp_1 \cache_data_B_reg[1][25]  ( .ip(n6207), .ck(clk), .q(
        \cache_data_B[1][25] ) );
  dp_1 \cache_data_B_reg[1][26]  ( .ip(n6206), .ck(clk), .q(
        \cache_data_B[1][26] ) );
  dp_1 \cache_data_B_reg[1][27]  ( .ip(n6205), .ck(clk), .q(
        \cache_data_B[1][27] ) );
  dp_1 \cache_data_B_reg[1][28]  ( .ip(n6204), .ck(clk), .q(
        \cache_data_B[1][28] ) );
  dp_1 \cache_data_B_reg[1][29]  ( .ip(n6203), .ck(clk), .q(
        \cache_data_B[1][29] ) );
  dp_1 \cache_data_B_reg[1][30]  ( .ip(n6202), .ck(clk), .q(
        \cache_data_B[1][30] ) );
  dp_1 \cache_data_B_reg[1][31]  ( .ip(n6201), .ck(clk), .q(
        \cache_data_B[1][31] ) );
  dp_1 \cache_data_B_reg[2][30]  ( .ip(n6104), .ck(clk), .q(
        \cache_data_B[2][30] ) );
  dp_1 \cache_data_B_reg[2][31]  ( .ip(n6103), .ck(clk), .q(
        \cache_data_B[2][31] ) );
  dp_1 \cache_data_B_reg[2][0]  ( .ip(n6102), .ck(clk), .q(
        \cache_data_B[2][0] ) );
  dp_1 \cache_data_B_reg[2][1]  ( .ip(n6101), .ck(clk), .q(
        \cache_data_B[2][1] ) );
  dp_1 \cache_data_B_reg[2][2]  ( .ip(n6100), .ck(clk), .q(
        \cache_data_B[2][2] ) );
  dp_1 \cache_data_B_reg[2][3]  ( .ip(n6099), .ck(clk), .q(
        \cache_data_B[2][3] ) );
  dp_1 \cache_data_B_reg[2][4]  ( .ip(n6098), .ck(clk), .q(
        \cache_data_B[2][4] ) );
  dp_1 \cache_data_B_reg[2][5]  ( .ip(n6097), .ck(clk), .q(
        \cache_data_B[2][5] ) );
  dp_1 \cache_data_B_reg[2][6]  ( .ip(n6096), .ck(clk), .q(
        \cache_data_B[2][6] ) );
  dp_1 \cache_data_B_reg[2][7]  ( .ip(n6095), .ck(clk), .q(
        \cache_data_B[2][7] ) );
  dp_1 \cache_data_B_reg[2][8]  ( .ip(n6094), .ck(clk), .q(
        \cache_data_B[2][8] ) );
  dp_1 \cache_data_B_reg[2][9]  ( .ip(n6093), .ck(clk), .q(
        \cache_data_B[2][9] ) );
  dp_1 \cache_data_B_reg[2][10]  ( .ip(n6092), .ck(clk), .q(
        \cache_data_B[2][10] ) );
  dp_1 \cache_data_B_reg[2][11]  ( .ip(n6091), .ck(clk), .q(
        \cache_data_B[2][11] ) );
  dp_1 \cache_data_B_reg[2][12]  ( .ip(n6090), .ck(clk), .q(
        \cache_data_B[2][12] ) );
  dp_1 \cache_data_B_reg[2][13]  ( .ip(n6089), .ck(clk), .q(
        \cache_data_B[2][13] ) );
  dp_1 \cache_data_B_reg[2][14]  ( .ip(n6088), .ck(clk), .q(
        \cache_data_B[2][14] ) );
  dp_1 \cache_data_B_reg[2][15]  ( .ip(n6087), .ck(clk), .q(
        \cache_data_B[2][15] ) );
  dp_1 \cache_data_B_reg[2][16]  ( .ip(n6086), .ck(clk), .q(
        \cache_data_B[2][16] ) );
  dp_1 \cache_data_B_reg[2][17]  ( .ip(n6085), .ck(clk), .q(
        \cache_data_B[2][17] ) );
  dp_1 \cache_data_B_reg[2][18]  ( .ip(n6084), .ck(clk), .q(
        \cache_data_B[2][18] ) );
  dp_1 \cache_data_B_reg[2][19]  ( .ip(n6083), .ck(clk), .q(
        \cache_data_B[2][19] ) );
  dp_1 \cache_data_B_reg[2][20]  ( .ip(n6082), .ck(clk), .q(
        \cache_data_B[2][20] ) );
  dp_1 \cache_data_B_reg[2][21]  ( .ip(n6081), .ck(clk), .q(
        \cache_data_B[2][21] ) );
  dp_1 \cache_data_B_reg[2][22]  ( .ip(n6080), .ck(clk), .q(
        \cache_data_B[2][22] ) );
  dp_1 \cache_data_B_reg[2][23]  ( .ip(n6079), .ck(clk), .q(
        \cache_data_B[2][23] ) );
  dp_1 \cache_data_B_reg[2][24]  ( .ip(n6078), .ck(clk), .q(
        \cache_data_B[2][24] ) );
  dp_1 \cache_data_B_reg[2][25]  ( .ip(n6077), .ck(clk), .q(
        \cache_data_B[2][25] ) );
  dp_1 \cache_data_B_reg[2][26]  ( .ip(n6076), .ck(clk), .q(
        \cache_data_B[2][26] ) );
  dp_1 \cache_data_B_reg[2][27]  ( .ip(n6075), .ck(clk), .q(
        \cache_data_B[2][27] ) );
  dp_1 \cache_data_B_reg[2][28]  ( .ip(n6074), .ck(clk), .q(
        \cache_data_B[2][28] ) );
  dp_1 \cache_data_B_reg[2][29]  ( .ip(n6073), .ck(clk), .q(
        \cache_data_B[2][29] ) );
  dp_1 \cache_data_B_reg[3][1]  ( .ip(n5976), .ck(clk), .q(
        \cache_data_B[3][1] ) );
  dp_1 \cache_data_B_reg[3][2]  ( .ip(n5975), .ck(clk), .q(
        \cache_data_B[3][2] ) );
  dp_1 \cache_data_B_reg[3][3]  ( .ip(n5974), .ck(clk), .q(
        \cache_data_B[3][3] ) );
  dp_1 \cache_data_B_reg[3][4]  ( .ip(n5973), .ck(clk), .q(
        \cache_data_B[3][4] ) );
  dp_1 \cache_data_B_reg[3][5]  ( .ip(n5972), .ck(clk), .q(
        \cache_data_B[3][5] ) );
  dp_1 \cache_data_B_reg[3][6]  ( .ip(n5971), .ck(clk), .q(
        \cache_data_B[3][6] ) );
  dp_1 \cache_data_B_reg[3][7]  ( .ip(n5970), .ck(clk), .q(
        \cache_data_B[3][7] ) );
  dp_1 \cache_data_B_reg[3][8]  ( .ip(n5969), .ck(clk), .q(
        \cache_data_B[3][8] ) );
  dp_1 \cache_data_B_reg[3][9]  ( .ip(n5968), .ck(clk), .q(
        \cache_data_B[3][9] ) );
  dp_1 \cache_data_B_reg[3][10]  ( .ip(n5967), .ck(clk), .q(
        \cache_data_B[3][10] ) );
  dp_1 \cache_data_B_reg[3][11]  ( .ip(n5966), .ck(clk), .q(
        \cache_data_B[3][11] ) );
  dp_1 \cache_data_B_reg[3][12]  ( .ip(n5965), .ck(clk), .q(
        \cache_data_B[3][12] ) );
  dp_1 \cache_data_B_reg[3][13]  ( .ip(n5964), .ck(clk), .q(
        \cache_data_B[3][13] ) );
  dp_1 \cache_data_B_reg[3][14]  ( .ip(n5963), .ck(clk), .q(
        \cache_data_B[3][14] ) );
  dp_1 \cache_data_B_reg[3][15]  ( .ip(n5962), .ck(clk), .q(
        \cache_data_B[3][15] ) );
  dp_1 \cache_data_B_reg[3][16]  ( .ip(n5961), .ck(clk), .q(
        \cache_data_B[3][16] ) );
  dp_1 \cache_data_B_reg[3][17]  ( .ip(n5960), .ck(clk), .q(
        \cache_data_B[3][17] ) );
  dp_1 \cache_data_B_reg[3][18]  ( .ip(n5959), .ck(clk), .q(
        \cache_data_B[3][18] ) );
  dp_1 \cache_data_B_reg[3][19]  ( .ip(n5958), .ck(clk), .q(
        \cache_data_B[3][19] ) );
  dp_1 \cache_data_B_reg[3][20]  ( .ip(n5957), .ck(clk), .q(
        \cache_data_B[3][20] ) );
  dp_1 \cache_data_B_reg[3][21]  ( .ip(n5956), .ck(clk), .q(
        \cache_data_B[3][21] ) );
  dp_1 \cache_data_B_reg[3][22]  ( .ip(n5955), .ck(clk), .q(
        \cache_data_B[3][22] ) );
  dp_1 \cache_data_B_reg[3][23]  ( .ip(n5954), .ck(clk), .q(
        \cache_data_B[3][23] ) );
  dp_1 \cache_data_B_reg[3][24]  ( .ip(n5953), .ck(clk), .q(
        \cache_data_B[3][24] ) );
  dp_1 \cache_data_B_reg[3][25]  ( .ip(n5952), .ck(clk), .q(
        \cache_data_B[3][25] ) );
  dp_1 \cache_data_B_reg[3][26]  ( .ip(n5951), .ck(clk), .q(
        \cache_data_B[3][26] ) );
  dp_1 \cache_data_B_reg[3][27]  ( .ip(n5950), .ck(clk), .q(
        \cache_data_B[3][27] ) );
  dp_1 \cache_data_B_reg[3][28]  ( .ip(n5949), .ck(clk), .q(
        \cache_data_B[3][28] ) );
  dp_1 \cache_data_B_reg[3][29]  ( .ip(n5948), .ck(clk), .q(
        \cache_data_B[3][29] ) );
  dp_1 \cache_data_B_reg[3][30]  ( .ip(n5947), .ck(clk), .q(
        \cache_data_B[3][30] ) );
  dp_1 \cache_data_B_reg[3][31]  ( .ip(n5946), .ck(clk), .q(
        \cache_data_B[3][31] ) );
  dp_1 \cache_data_B_reg[3][0]  ( .ip(n5945), .ck(clk), .q(
        \cache_data_B[3][0] ) );
  dp_1 \cache_data_B_reg[4][0]  ( .ip(n5848), .ck(clk), .q(
        \cache_data_B[4][0] ) );
  dp_1 \cache_data_B_reg[4][1]  ( .ip(n5847), .ck(clk), .q(
        \cache_data_B[4][1] ) );
  dp_1 \cache_data_B_reg[4][2]  ( .ip(n5846), .ck(clk), .q(
        \cache_data_B[4][2] ) );
  dp_1 \cache_data_B_reg[4][3]  ( .ip(n5845), .ck(clk), .q(
        \cache_data_B[4][3] ) );
  dp_1 \cache_data_B_reg[4][4]  ( .ip(n5844), .ck(clk), .q(
        \cache_data_B[4][4] ) );
  dp_1 \cache_data_B_reg[4][5]  ( .ip(n5843), .ck(clk), .q(
        \cache_data_B[4][5] ) );
  dp_1 \cache_data_B_reg[4][6]  ( .ip(n5842), .ck(clk), .q(
        \cache_data_B[4][6] ) );
  dp_1 \cache_data_B_reg[4][7]  ( .ip(n5841), .ck(clk), .q(
        \cache_data_B[4][7] ) );
  dp_1 \cache_data_B_reg[4][8]  ( .ip(n5840), .ck(clk), .q(
        \cache_data_B[4][8] ) );
  dp_1 \cache_data_B_reg[4][9]  ( .ip(n5839), .ck(clk), .q(
        \cache_data_B[4][9] ) );
  dp_1 \cache_data_B_reg[4][10]  ( .ip(n5838), .ck(clk), .q(
        \cache_data_B[4][10] ) );
  dp_1 \cache_data_B_reg[4][11]  ( .ip(n5837), .ck(clk), .q(
        \cache_data_B[4][11] ) );
  dp_1 \cache_data_B_reg[4][12]  ( .ip(n5836), .ck(clk), .q(
        \cache_data_B[4][12] ) );
  dp_1 \cache_data_B_reg[4][13]  ( .ip(n5835), .ck(clk), .q(
        \cache_data_B[4][13] ) );
  dp_1 \cache_data_B_reg[4][14]  ( .ip(n5834), .ck(clk), .q(
        \cache_data_B[4][14] ) );
  dp_1 \cache_data_B_reg[4][15]  ( .ip(n5833), .ck(clk), .q(
        \cache_data_B[4][15] ) );
  dp_1 \cache_data_B_reg[4][16]  ( .ip(n5832), .ck(clk), .q(
        \cache_data_B[4][16] ) );
  dp_1 \cache_data_B_reg[4][17]  ( .ip(n5831), .ck(clk), .q(
        \cache_data_B[4][17] ) );
  dp_1 \cache_data_B_reg[4][18]  ( .ip(n5830), .ck(clk), .q(
        \cache_data_B[4][18] ) );
  dp_1 \cache_data_B_reg[4][19]  ( .ip(n5829), .ck(clk), .q(
        \cache_data_B[4][19] ) );
  dp_1 \cache_data_B_reg[4][20]  ( .ip(n5828), .ck(clk), .q(
        \cache_data_B[4][20] ) );
  dp_1 \cache_data_B_reg[4][21]  ( .ip(n5827), .ck(clk), .q(
        \cache_data_B[4][21] ) );
  dp_1 \cache_data_B_reg[4][22]  ( .ip(n5826), .ck(clk), .q(
        \cache_data_B[4][22] ) );
  dp_1 \cache_data_B_reg[4][23]  ( .ip(n5825), .ck(clk), .q(
        \cache_data_B[4][23] ) );
  dp_1 \cache_data_B_reg[4][24]  ( .ip(n5824), .ck(clk), .q(
        \cache_data_B[4][24] ) );
  dp_1 \cache_data_B_reg[4][25]  ( .ip(n5823), .ck(clk), .q(
        \cache_data_B[4][25] ) );
  dp_1 \cache_data_B_reg[4][26]  ( .ip(n5822), .ck(clk), .q(
        \cache_data_B[4][26] ) );
  dp_1 \cache_data_B_reg[4][27]  ( .ip(n5821), .ck(clk), .q(
        \cache_data_B[4][27] ) );
  dp_1 \cache_data_B_reg[4][28]  ( .ip(n5820), .ck(clk), .q(
        \cache_data_B[4][28] ) );
  dp_1 \cache_data_B_reg[4][29]  ( .ip(n5819), .ck(clk), .q(
        \cache_data_B[4][29] ) );
  dp_1 \cache_data_B_reg[4][30]  ( .ip(n5818), .ck(clk), .q(
        \cache_data_B[4][30] ) );
  dp_1 \cache_data_B_reg[4][31]  ( .ip(n5817), .ck(clk), .q(
        \cache_data_B[4][31] ) );
  dp_1 \cache_data_B_reg[5][0]  ( .ip(n5720), .ck(clk), .q(
        \cache_data_B[5][0] ) );
  dp_1 \cache_data_B_reg[5][1]  ( .ip(n5719), .ck(clk), .q(
        \cache_data_B[5][1] ) );
  dp_1 \cache_data_B_reg[5][2]  ( .ip(n5718), .ck(clk), .q(
        \cache_data_B[5][2] ) );
  dp_1 \cache_data_B_reg[5][3]  ( .ip(n5717), .ck(clk), .q(
        \cache_data_B[5][3] ) );
  dp_1 \cache_data_B_reg[5][4]  ( .ip(n5716), .ck(clk), .q(
        \cache_data_B[5][4] ) );
  dp_1 \cache_data_B_reg[5][5]  ( .ip(n5715), .ck(clk), .q(
        \cache_data_B[5][5] ) );
  dp_1 \cache_data_B_reg[5][6]  ( .ip(n5714), .ck(clk), .q(
        \cache_data_B[5][6] ) );
  dp_1 \cache_data_B_reg[5][7]  ( .ip(n5713), .ck(clk), .q(
        \cache_data_B[5][7] ) );
  dp_1 \cache_data_B_reg[5][8]  ( .ip(n5712), .ck(clk), .q(
        \cache_data_B[5][8] ) );
  dp_1 \cache_data_B_reg[5][9]  ( .ip(n5711), .ck(clk), .q(
        \cache_data_B[5][9] ) );
  dp_1 \cache_data_B_reg[5][10]  ( .ip(n5710), .ck(clk), .q(
        \cache_data_B[5][10] ) );
  dp_1 \cache_data_B_reg[5][11]  ( .ip(n5709), .ck(clk), .q(
        \cache_data_B[5][11] ) );
  dp_1 \cache_data_B_reg[5][12]  ( .ip(n5708), .ck(clk), .q(
        \cache_data_B[5][12] ) );
  dp_1 \cache_data_B_reg[5][13]  ( .ip(n5707), .ck(clk), .q(
        \cache_data_B[5][13] ) );
  dp_1 \cache_data_B_reg[5][14]  ( .ip(n5706), .ck(clk), .q(
        \cache_data_B[5][14] ) );
  dp_1 \cache_data_B_reg[5][15]  ( .ip(n5705), .ck(clk), .q(
        \cache_data_B[5][15] ) );
  dp_1 \cache_data_B_reg[5][16]  ( .ip(n5704), .ck(clk), .q(
        \cache_data_B[5][16] ) );
  dp_1 \cache_data_B_reg[5][17]  ( .ip(n5703), .ck(clk), .q(
        \cache_data_B[5][17] ) );
  dp_1 \cache_data_B_reg[5][18]  ( .ip(n5702), .ck(clk), .q(
        \cache_data_B[5][18] ) );
  dp_1 \cache_data_B_reg[5][19]  ( .ip(n5701), .ck(clk), .q(
        \cache_data_B[5][19] ) );
  dp_1 \cache_data_B_reg[5][20]  ( .ip(n5700), .ck(clk), .q(
        \cache_data_B[5][20] ) );
  dp_1 \cache_data_B_reg[5][21]  ( .ip(n5699), .ck(clk), .q(
        \cache_data_B[5][21] ) );
  dp_1 \cache_data_B_reg[5][22]  ( .ip(n5698), .ck(clk), .q(
        \cache_data_B[5][22] ) );
  dp_1 \cache_data_B_reg[5][23]  ( .ip(n5697), .ck(clk), .q(
        \cache_data_B[5][23] ) );
  dp_1 \cache_data_B_reg[5][24]  ( .ip(n5696), .ck(clk), .q(
        \cache_data_B[5][24] ) );
  dp_1 \cache_data_B_reg[5][25]  ( .ip(n5695), .ck(clk), .q(
        \cache_data_B[5][25] ) );
  dp_1 \cache_data_B_reg[5][26]  ( .ip(n5694), .ck(clk), .q(
        \cache_data_B[5][26] ) );
  dp_1 \cache_data_B_reg[5][27]  ( .ip(n5693), .ck(clk), .q(
        \cache_data_B[5][27] ) );
  dp_1 \cache_data_B_reg[5][28]  ( .ip(n5692), .ck(clk), .q(
        \cache_data_B[5][28] ) );
  dp_1 \cache_data_B_reg[5][29]  ( .ip(n5691), .ck(clk), .q(
        \cache_data_B[5][29] ) );
  dp_1 \cache_data_B_reg[5][30]  ( .ip(n5690), .ck(clk), .q(
        \cache_data_B[5][30] ) );
  dp_1 \cache_data_B_reg[5][31]  ( .ip(n5689), .ck(clk), .q(
        \cache_data_B[5][31] ) );
  dp_1 \cache_data_B_reg[6][13]  ( .ip(n5592), .ck(clk), .q(
        \cache_data_B[6][13] ) );
  dp_1 \cache_data_B_reg[6][14]  ( .ip(n5591), .ck(clk), .q(
        \cache_data_B[6][14] ) );
  dp_1 \cache_data_B_reg[6][15]  ( .ip(n5590), .ck(clk), .q(
        \cache_data_B[6][15] ) );
  dp_1 \cache_data_B_reg[6][16]  ( .ip(n5589), .ck(clk), .q(
        \cache_data_B[6][16] ) );
  dp_1 \cache_data_B_reg[6][17]  ( .ip(n5588), .ck(clk), .q(
        \cache_data_B[6][17] ) );
  dp_1 \cache_data_B_reg[6][18]  ( .ip(n5587), .ck(clk), .q(
        \cache_data_B[6][18] ) );
  dp_1 \cache_data_B_reg[6][19]  ( .ip(n5586), .ck(clk), .q(
        \cache_data_B[6][19] ) );
  dp_1 \cache_data_B_reg[6][20]  ( .ip(n5585), .ck(clk), .q(
        \cache_data_B[6][20] ) );
  dp_1 \cache_data_B_reg[6][21]  ( .ip(n5584), .ck(clk), .q(
        \cache_data_B[6][21] ) );
  dp_1 \cache_data_B_reg[6][22]  ( .ip(n5583), .ck(clk), .q(
        \cache_data_B[6][22] ) );
  dp_1 \cache_data_B_reg[6][23]  ( .ip(n5582), .ck(clk), .q(
        \cache_data_B[6][23] ) );
  dp_1 \cache_data_B_reg[6][24]  ( .ip(n5581), .ck(clk), .q(
        \cache_data_B[6][24] ) );
  dp_1 \cache_data_B_reg[6][25]  ( .ip(n5580), .ck(clk), .q(
        \cache_data_B[6][25] ) );
  dp_1 \cache_data_B_reg[6][26]  ( .ip(n5579), .ck(clk), .q(
        \cache_data_B[6][26] ) );
  dp_1 \cache_data_B_reg[6][27]  ( .ip(n5578), .ck(clk), .q(
        \cache_data_B[6][27] ) );
  dp_1 \cache_data_B_reg[6][28]  ( .ip(n5577), .ck(clk), .q(
        \cache_data_B[6][28] ) );
  dp_1 \cache_data_B_reg[6][29]  ( .ip(n5576), .ck(clk), .q(
        \cache_data_B[6][29] ) );
  dp_1 \cache_data_B_reg[6][30]  ( .ip(n5575), .ck(clk), .q(
        \cache_data_B[6][30] ) );
  dp_1 \cache_data_B_reg[6][31]  ( .ip(n5574), .ck(clk), .q(
        \cache_data_B[6][31] ) );
  dp_1 \cache_data_B_reg[6][0]  ( .ip(n5573), .ck(clk), .q(
        \cache_data_B[6][0] ) );
  dp_1 \cache_data_B_reg[6][1]  ( .ip(n5572), .ck(clk), .q(
        \cache_data_B[6][1] ) );
  dp_1 \cache_data_B_reg[6][2]  ( .ip(n5571), .ck(clk), .q(
        \cache_data_B[6][2] ) );
  dp_1 \cache_data_B_reg[6][3]  ( .ip(n5570), .ck(clk), .q(
        \cache_data_B[6][3] ) );
  dp_1 \cache_data_B_reg[6][4]  ( .ip(n5569), .ck(clk), .q(
        \cache_data_B[6][4] ) );
  dp_1 \cache_data_B_reg[6][5]  ( .ip(n5568), .ck(clk), .q(
        \cache_data_B[6][5] ) );
  dp_1 \cache_data_B_reg[6][6]  ( .ip(n5567), .ck(clk), .q(
        \cache_data_B[6][6] ) );
  dp_1 \cache_data_B_reg[6][7]  ( .ip(n5566), .ck(clk), .q(
        \cache_data_B[6][7] ) );
  dp_1 \cache_data_B_reg[6][8]  ( .ip(n5565), .ck(clk), .q(
        \cache_data_B[6][8] ) );
  dp_1 \cache_data_B_reg[6][9]  ( .ip(n5564), .ck(clk), .q(
        \cache_data_B[6][9] ) );
  dp_1 \cache_data_B_reg[6][10]  ( .ip(n5563), .ck(clk), .q(
        \cache_data_B[6][10] ) );
  dp_1 \cache_data_B_reg[6][11]  ( .ip(n5562), .ck(clk), .q(
        \cache_data_B[6][11] ) );
  dp_1 \cache_data_B_reg[6][12]  ( .ip(n5561), .ck(clk), .q(
        \cache_data_B[6][12] ) );
  dp_1 \cache_data_B_reg[7][0]  ( .ip(n5464), .ck(clk), .q(
        \cache_data_B[7][0] ) );
  dp_1 \cache_data_B_reg[7][1]  ( .ip(n5463), .ck(clk), .q(
        \cache_data_B[7][1] ) );
  dp_1 \cache_data_B_reg[7][2]  ( .ip(n5462), .ck(clk), .q(
        \cache_data_B[7][2] ) );
  dp_1 \cache_data_B_reg[7][3]  ( .ip(n5461), .ck(clk), .q(
        \cache_data_B[7][3] ) );
  dp_1 \cache_data_B_reg[7][4]  ( .ip(n5460), .ck(clk), .q(
        \cache_data_B[7][4] ) );
  dp_1 \cache_data_B_reg[7][5]  ( .ip(n5459), .ck(clk), .q(
        \cache_data_B[7][5] ) );
  dp_1 \cache_data_B_reg[7][6]  ( .ip(n5458), .ck(clk), .q(
        \cache_data_B[7][6] ) );
  dp_1 \cache_data_B_reg[7][7]  ( .ip(n5457), .ck(clk), .q(
        \cache_data_B[7][7] ) );
  dp_1 \cache_data_B_reg[7][8]  ( .ip(n5456), .ck(clk), .q(
        \cache_data_B[7][8] ) );
  dp_1 \cache_data_B_reg[7][9]  ( .ip(n5455), .ck(clk), .q(
        \cache_data_B[7][9] ) );
  dp_1 \cache_data_B_reg[7][10]  ( .ip(n5454), .ck(clk), .q(
        \cache_data_B[7][10] ) );
  dp_1 \cache_data_B_reg[7][11]  ( .ip(n5453), .ck(clk), .q(
        \cache_data_B[7][11] ) );
  dp_1 \cache_data_B_reg[7][12]  ( .ip(n5452), .ck(clk), .q(
        \cache_data_B[7][12] ) );
  dp_1 \cache_data_B_reg[7][13]  ( .ip(n5451), .ck(clk), .q(
        \cache_data_B[7][13] ) );
  dp_1 \cache_data_B_reg[7][14]  ( .ip(n5450), .ck(clk), .q(
        \cache_data_B[7][14] ) );
  dp_1 \cache_data_B_reg[7][15]  ( .ip(n5449), .ck(clk), .q(
        \cache_data_B[7][15] ) );
  dp_1 \cache_data_B_reg[7][16]  ( .ip(n5448), .ck(clk), .q(
        \cache_data_B[7][16] ) );
  dp_1 \cache_data_B_reg[7][17]  ( .ip(n5447), .ck(clk), .q(
        \cache_data_B[7][17] ) );
  dp_1 \cache_data_B_reg[7][18]  ( .ip(n5446), .ck(clk), .q(
        \cache_data_B[7][18] ) );
  dp_1 \cache_data_B_reg[7][19]  ( .ip(n5445), .ck(clk), .q(
        \cache_data_B[7][19] ) );
  dp_1 \cache_data_B_reg[7][20]  ( .ip(n5444), .ck(clk), .q(
        \cache_data_B[7][20] ) );
  dp_1 \cache_data_B_reg[7][21]  ( .ip(n5443), .ck(clk), .q(
        \cache_data_B[7][21] ) );
  dp_1 \cache_data_B_reg[7][22]  ( .ip(n5442), .ck(clk), .q(
        \cache_data_B[7][22] ) );
  dp_1 \cache_data_B_reg[7][23]  ( .ip(n5441), .ck(clk), .q(
        \cache_data_B[7][23] ) );
  dp_1 \cache_data_B_reg[7][24]  ( .ip(n5440), .ck(clk), .q(
        \cache_data_B[7][24] ) );
  dp_1 \cache_data_B_reg[7][25]  ( .ip(n5439), .ck(clk), .q(
        \cache_data_B[7][25] ) );
  dp_1 \cache_data_B_reg[7][26]  ( .ip(n5438), .ck(clk), .q(
        \cache_data_B[7][26] ) );
  dp_1 \cache_data_B_reg[7][27]  ( .ip(n5437), .ck(clk), .q(
        \cache_data_B[7][27] ) );
  dp_1 \cache_data_B_reg[7][28]  ( .ip(n5436), .ck(clk), .q(
        \cache_data_B[7][28] ) );
  dp_1 \cache_data_B_reg[7][29]  ( .ip(n5435), .ck(clk), .q(
        \cache_data_B[7][29] ) );
  dp_1 \cache_data_B_reg[7][30]  ( .ip(n5434), .ck(clk), .q(
        \cache_data_B[7][30] ) );
  dp_1 \cache_data_B_reg[7][31]  ( .ip(n5433), .ck(clk), .q(
        \cache_data_B[7][31] ) );
  dp_1 \cache_data_B_reg[0][32]  ( .ip(n6328), .ck(clk), .q(
        \cache_data_B[0][32] ) );
  dp_1 \cache_data_B_reg[0][33]  ( .ip(n6327), .ck(clk), .q(
        \cache_data_B[0][33] ) );
  dp_1 \cache_data_B_reg[0][34]  ( .ip(n6326), .ck(clk), .q(
        \cache_data_B[0][34] ) );
  dp_1 \cache_data_B_reg[0][35]  ( .ip(n6325), .ck(clk), .q(
        \cache_data_B[0][35] ) );
  dp_1 \cache_data_B_reg[0][36]  ( .ip(n6324), .ck(clk), .q(
        \cache_data_B[0][36] ) );
  dp_1 \cache_data_B_reg[0][37]  ( .ip(n6323), .ck(clk), .q(
        \cache_data_B[0][37] ) );
  dp_1 \cache_data_B_reg[0][38]  ( .ip(n6322), .ck(clk), .q(
        \cache_data_B[0][38] ) );
  dp_1 \cache_data_B_reg[0][39]  ( .ip(n6321), .ck(clk), .q(
        \cache_data_B[0][39] ) );
  dp_1 \cache_data_B_reg[0][40]  ( .ip(n6320), .ck(clk), .q(
        \cache_data_B[0][40] ) );
  dp_1 \cache_data_B_reg[0][41]  ( .ip(n6319), .ck(clk), .q(
        \cache_data_B[0][41] ) );
  dp_1 \cache_data_B_reg[0][42]  ( .ip(n6318), .ck(clk), .q(
        \cache_data_B[0][42] ) );
  dp_1 \cache_data_B_reg[0][43]  ( .ip(n6317), .ck(clk), .q(
        \cache_data_B[0][43] ) );
  dp_1 \cache_data_B_reg[0][44]  ( .ip(n6316), .ck(clk), .q(
        \cache_data_B[0][44] ) );
  dp_1 \cache_data_B_reg[0][45]  ( .ip(n6315), .ck(clk), .q(
        \cache_data_B[0][45] ) );
  dp_1 \cache_data_B_reg[0][46]  ( .ip(n6314), .ck(clk), .q(
        \cache_data_B[0][46] ) );
  dp_1 \cache_data_B_reg[0][47]  ( .ip(n6313), .ck(clk), .q(
        \cache_data_B[0][47] ) );
  dp_1 \cache_data_B_reg[0][48]  ( .ip(n6312), .ck(clk), .q(
        \cache_data_B[0][48] ) );
  dp_1 \cache_data_B_reg[0][49]  ( .ip(n6311), .ck(clk), .q(
        \cache_data_B[0][49] ) );
  dp_1 \cache_data_B_reg[0][50]  ( .ip(n6310), .ck(clk), .q(
        \cache_data_B[0][50] ) );
  dp_1 \cache_data_B_reg[0][51]  ( .ip(n6309), .ck(clk), .q(
        \cache_data_B[0][51] ) );
  dp_1 \cache_data_B_reg[0][52]  ( .ip(n6308), .ck(clk), .q(
        \cache_data_B[0][52] ) );
  dp_1 \cache_data_B_reg[0][53]  ( .ip(n6307), .ck(clk), .q(
        \cache_data_B[0][53] ) );
  dp_1 \cache_data_B_reg[0][54]  ( .ip(n6306), .ck(clk), .q(
        \cache_data_B[0][54] ) );
  dp_1 \cache_data_B_reg[0][55]  ( .ip(n6305), .ck(clk), .q(
        \cache_data_B[0][55] ) );
  dp_1 \cache_data_B_reg[0][56]  ( .ip(n6304), .ck(clk), .q(
        \cache_data_B[0][56] ) );
  dp_1 \cache_data_B_reg[0][57]  ( .ip(n6303), .ck(clk), .q(
        \cache_data_B[0][57] ) );
  dp_1 \cache_data_B_reg[0][58]  ( .ip(n6302), .ck(clk), .q(
        \cache_data_B[0][58] ) );
  dp_1 \cache_data_B_reg[0][59]  ( .ip(n6301), .ck(clk), .q(
        \cache_data_B[0][59] ) );
  dp_1 \cache_data_B_reg[0][60]  ( .ip(n6300), .ck(clk), .q(
        \cache_data_B[0][60] ) );
  dp_1 \cache_data_B_reg[0][61]  ( .ip(n6299), .ck(clk), .q(
        \cache_data_B[0][61] ) );
  dp_1 \cache_data_B_reg[0][62]  ( .ip(n6298), .ck(clk), .q(
        \cache_data_B[0][62] ) );
  dp_1 \cache_data_B_reg[0][63]  ( .ip(n6297), .ck(clk), .q(
        \cache_data_B[0][63] ) );
  dp_1 \cache_data_B_reg[1][59]  ( .ip(n6200), .ck(clk), .q(
        \cache_data_B[1][59] ) );
  dp_1 \cache_data_B_reg[1][60]  ( .ip(n6199), .ck(clk), .q(
        \cache_data_B[1][60] ) );
  dp_1 \cache_data_B_reg[1][61]  ( .ip(n6198), .ck(clk), .q(
        \cache_data_B[1][61] ) );
  dp_1 \cache_data_B_reg[1][62]  ( .ip(n6197), .ck(clk), .q(
        \cache_data_B[1][62] ) );
  dp_1 \cache_data_B_reg[1][63]  ( .ip(n6196), .ck(clk), .q(
        \cache_data_B[1][63] ) );
  dp_1 \cache_data_B_reg[1][32]  ( .ip(n6195), .ck(clk), .q(
        \cache_data_B[1][32] ) );
  dp_1 \cache_data_B_reg[1][33]  ( .ip(n6194), .ck(clk), .q(
        \cache_data_B[1][33] ) );
  dp_1 \cache_data_B_reg[1][34]  ( .ip(n6193), .ck(clk), .q(
        \cache_data_B[1][34] ) );
  dp_1 \cache_data_B_reg[1][35]  ( .ip(n6192), .ck(clk), .q(
        \cache_data_B[1][35] ) );
  dp_1 \cache_data_B_reg[1][36]  ( .ip(n6191), .ck(clk), .q(
        \cache_data_B[1][36] ) );
  dp_1 \cache_data_B_reg[1][37]  ( .ip(n6190), .ck(clk), .q(
        \cache_data_B[1][37] ) );
  dp_1 \cache_data_B_reg[1][38]  ( .ip(n6189), .ck(clk), .q(
        \cache_data_B[1][38] ) );
  dp_1 \cache_data_B_reg[1][39]  ( .ip(n6188), .ck(clk), .q(
        \cache_data_B[1][39] ) );
  dp_1 \cache_data_B_reg[1][40]  ( .ip(n6187), .ck(clk), .q(
        \cache_data_B[1][40] ) );
  dp_1 \cache_data_B_reg[1][41]  ( .ip(n6186), .ck(clk), .q(
        \cache_data_B[1][41] ) );
  dp_1 \cache_data_B_reg[1][42]  ( .ip(n6185), .ck(clk), .q(
        \cache_data_B[1][42] ) );
  dp_1 \cache_data_B_reg[1][43]  ( .ip(n6184), .ck(clk), .q(
        \cache_data_B[1][43] ) );
  dp_1 \cache_data_B_reg[1][44]  ( .ip(n6183), .ck(clk), .q(
        \cache_data_B[1][44] ) );
  dp_1 \cache_data_B_reg[1][45]  ( .ip(n6182), .ck(clk), .q(
        \cache_data_B[1][45] ) );
  dp_1 \cache_data_B_reg[1][46]  ( .ip(n6181), .ck(clk), .q(
        \cache_data_B[1][46] ) );
  dp_1 \cache_data_B_reg[1][47]  ( .ip(n6180), .ck(clk), .q(
        \cache_data_B[1][47] ) );
  dp_1 \cache_data_B_reg[1][48]  ( .ip(n6179), .ck(clk), .q(
        \cache_data_B[1][48] ) );
  dp_1 \cache_data_B_reg[1][49]  ( .ip(n6178), .ck(clk), .q(
        \cache_data_B[1][49] ) );
  dp_1 \cache_data_B_reg[1][50]  ( .ip(n6177), .ck(clk), .q(
        \cache_data_B[1][50] ) );
  dp_1 \cache_data_B_reg[1][51]  ( .ip(n6176), .ck(clk), .q(
        \cache_data_B[1][51] ) );
  dp_1 \cache_data_B_reg[1][52]  ( .ip(n6175), .ck(clk), .q(
        \cache_data_B[1][52] ) );
  dp_1 \cache_data_B_reg[1][53]  ( .ip(n6174), .ck(clk), .q(
        \cache_data_B[1][53] ) );
  dp_1 \cache_data_B_reg[1][54]  ( .ip(n6173), .ck(clk), .q(
        \cache_data_B[1][54] ) );
  dp_1 \cache_data_B_reg[1][55]  ( .ip(n6172), .ck(clk), .q(
        \cache_data_B[1][55] ) );
  dp_1 \cache_data_B_reg[1][56]  ( .ip(n6171), .ck(clk), .q(
        \cache_data_B[1][56] ) );
  dp_1 \cache_data_B_reg[1][57]  ( .ip(n6170), .ck(clk), .q(
        \cache_data_B[1][57] ) );
  dp_1 \cache_data_B_reg[1][58]  ( .ip(n6169), .ck(clk), .q(
        \cache_data_B[1][58] ) );
  dp_1 \cache_data_B_reg[2][32]  ( .ip(n6072), .ck(clk), .q(
        \cache_data_B[2][32] ) );
  dp_1 \cache_data_B_reg[2][33]  ( .ip(n6071), .ck(clk), .q(
        \cache_data_B[2][33] ) );
  dp_1 \cache_data_B_reg[2][34]  ( .ip(n6070), .ck(clk), .q(
        \cache_data_B[2][34] ) );
  dp_1 \cache_data_B_reg[2][35]  ( .ip(n6069), .ck(clk), .q(
        \cache_data_B[2][35] ) );
  dp_1 \cache_data_B_reg[2][36]  ( .ip(n6068), .ck(clk), .q(
        \cache_data_B[2][36] ) );
  dp_1 \cache_data_B_reg[2][37]  ( .ip(n6067), .ck(clk), .q(
        \cache_data_B[2][37] ) );
  dp_1 \cache_data_B_reg[2][38]  ( .ip(n6066), .ck(clk), .q(
        \cache_data_B[2][38] ) );
  dp_1 \cache_data_B_reg[2][39]  ( .ip(n6065), .ck(clk), .q(
        \cache_data_B[2][39] ) );
  dp_1 \cache_data_B_reg[2][40]  ( .ip(n6064), .ck(clk), .q(
        \cache_data_B[2][40] ) );
  dp_1 \cache_data_B_reg[2][41]  ( .ip(n6063), .ck(clk), .q(
        \cache_data_B[2][41] ) );
  dp_1 \cache_data_B_reg[2][42]  ( .ip(n6062), .ck(clk), .q(
        \cache_data_B[2][42] ) );
  dp_1 \cache_data_B_reg[2][43]  ( .ip(n6061), .ck(clk), .q(
        \cache_data_B[2][43] ) );
  dp_1 \cache_data_B_reg[2][44]  ( .ip(n6060), .ck(clk), .q(
        \cache_data_B[2][44] ) );
  dp_1 \cache_data_B_reg[2][45]  ( .ip(n6059), .ck(clk), .q(
        \cache_data_B[2][45] ) );
  dp_1 \cache_data_B_reg[2][46]  ( .ip(n6058), .ck(clk), .q(
        \cache_data_B[2][46] ) );
  dp_1 \cache_data_B_reg[2][47]  ( .ip(n6057), .ck(clk), .q(
        \cache_data_B[2][47] ) );
  dp_1 \cache_data_B_reg[2][48]  ( .ip(n6056), .ck(clk), .q(
        \cache_data_B[2][48] ) );
  dp_1 \cache_data_B_reg[2][49]  ( .ip(n6055), .ck(clk), .q(
        \cache_data_B[2][49] ) );
  dp_1 \cache_data_B_reg[2][50]  ( .ip(n6054), .ck(clk), .q(
        \cache_data_B[2][50] ) );
  dp_1 \cache_data_B_reg[2][51]  ( .ip(n6053), .ck(clk), .q(
        \cache_data_B[2][51] ) );
  dp_1 \cache_data_B_reg[2][52]  ( .ip(n6052), .ck(clk), .q(
        \cache_data_B[2][52] ) );
  dp_1 \cache_data_B_reg[2][53]  ( .ip(n6051), .ck(clk), .q(
        \cache_data_B[2][53] ) );
  dp_1 \cache_data_B_reg[2][54]  ( .ip(n6050), .ck(clk), .q(
        \cache_data_B[2][54] ) );
  dp_1 \cache_data_B_reg[2][55]  ( .ip(n6049), .ck(clk), .q(
        \cache_data_B[2][55] ) );
  dp_1 \cache_data_B_reg[2][56]  ( .ip(n6048), .ck(clk), .q(
        \cache_data_B[2][56] ) );
  dp_1 \cache_data_B_reg[2][57]  ( .ip(n6047), .ck(clk), .q(
        \cache_data_B[2][57] ) );
  dp_1 \cache_data_B_reg[2][58]  ( .ip(n6046), .ck(clk), .q(
        \cache_data_B[2][58] ) );
  dp_1 \cache_data_B_reg[2][59]  ( .ip(n6045), .ck(clk), .q(
        \cache_data_B[2][59] ) );
  dp_1 \cache_data_B_reg[2][60]  ( .ip(n6044), .ck(clk), .q(
        \cache_data_B[2][60] ) );
  dp_1 \cache_data_B_reg[2][61]  ( .ip(n6043), .ck(clk), .q(
        \cache_data_B[2][61] ) );
  dp_1 \cache_data_B_reg[2][62]  ( .ip(n6042), .ck(clk), .q(
        \cache_data_B[2][62] ) );
  dp_1 \cache_data_B_reg[2][63]  ( .ip(n6041), .ck(clk), .q(
        \cache_data_B[2][63] ) );
  dp_1 \cache_data_B_reg[3][32]  ( .ip(n5944), .ck(clk), .q(
        \cache_data_B[3][32] ) );
  dp_1 \cache_data_B_reg[3][33]  ( .ip(n5943), .ck(clk), .q(
        \cache_data_B[3][33] ) );
  dp_1 \cache_data_B_reg[3][34]  ( .ip(n5942), .ck(clk), .q(
        \cache_data_B[3][34] ) );
  dp_1 \cache_data_B_reg[3][35]  ( .ip(n5941), .ck(clk), .q(
        \cache_data_B[3][35] ) );
  dp_1 \cache_data_B_reg[3][36]  ( .ip(n5940), .ck(clk), .q(
        \cache_data_B[3][36] ) );
  dp_1 \cache_data_B_reg[3][37]  ( .ip(n5939), .ck(clk), .q(
        \cache_data_B[3][37] ) );
  dp_1 \cache_data_B_reg[3][38]  ( .ip(n5938), .ck(clk), .q(
        \cache_data_B[3][38] ) );
  dp_1 \cache_data_B_reg[3][39]  ( .ip(n5937), .ck(clk), .q(
        \cache_data_B[3][39] ) );
  dp_1 \cache_data_B_reg[3][40]  ( .ip(n5936), .ck(clk), .q(
        \cache_data_B[3][40] ) );
  dp_1 \cache_data_B_reg[3][41]  ( .ip(n5935), .ck(clk), .q(
        \cache_data_B[3][41] ) );
  dp_1 \cache_data_B_reg[3][42]  ( .ip(n5934), .ck(clk), .q(
        \cache_data_B[3][42] ) );
  dp_1 \cache_data_B_reg[3][43]  ( .ip(n5933), .ck(clk), .q(
        \cache_data_B[3][43] ) );
  dp_1 \cache_data_B_reg[3][44]  ( .ip(n5932), .ck(clk), .q(
        \cache_data_B[3][44] ) );
  dp_1 \cache_data_B_reg[3][45]  ( .ip(n5931), .ck(clk), .q(
        \cache_data_B[3][45] ) );
  dp_1 \cache_data_B_reg[3][46]  ( .ip(n5930), .ck(clk), .q(
        \cache_data_B[3][46] ) );
  dp_1 \cache_data_B_reg[3][47]  ( .ip(n5929), .ck(clk), .q(
        \cache_data_B[3][47] ) );
  dp_1 \cache_data_B_reg[3][48]  ( .ip(n5928), .ck(clk), .q(
        \cache_data_B[3][48] ) );
  dp_1 \cache_data_B_reg[3][49]  ( .ip(n5927), .ck(clk), .q(
        \cache_data_B[3][49] ) );
  dp_1 \cache_data_B_reg[3][50]  ( .ip(n5926), .ck(clk), .q(
        \cache_data_B[3][50] ) );
  dp_1 \cache_data_B_reg[3][51]  ( .ip(n5925), .ck(clk), .q(
        \cache_data_B[3][51] ) );
  dp_1 \cache_data_B_reg[3][52]  ( .ip(n5924), .ck(clk), .q(
        \cache_data_B[3][52] ) );
  dp_1 \cache_data_B_reg[3][53]  ( .ip(n5923), .ck(clk), .q(
        \cache_data_B[3][53] ) );
  dp_1 \cache_data_B_reg[3][54]  ( .ip(n5922), .ck(clk), .q(
        \cache_data_B[3][54] ) );
  dp_1 \cache_data_B_reg[3][55]  ( .ip(n5921), .ck(clk), .q(
        \cache_data_B[3][55] ) );
  dp_1 \cache_data_B_reg[3][56]  ( .ip(n5920), .ck(clk), .q(
        \cache_data_B[3][56] ) );
  dp_1 \cache_data_B_reg[3][57]  ( .ip(n5919), .ck(clk), .q(
        \cache_data_B[3][57] ) );
  dp_1 \cache_data_B_reg[3][58]  ( .ip(n5918), .ck(clk), .q(
        \cache_data_B[3][58] ) );
  dp_1 \cache_data_B_reg[3][59]  ( .ip(n5917), .ck(clk), .q(
        \cache_data_B[3][59] ) );
  dp_1 \cache_data_B_reg[3][60]  ( .ip(n5916), .ck(clk), .q(
        \cache_data_B[3][60] ) );
  dp_1 \cache_data_B_reg[3][61]  ( .ip(n5915), .ck(clk), .q(
        \cache_data_B[3][61] ) );
  dp_1 \cache_data_B_reg[3][62]  ( .ip(n5914), .ck(clk), .q(
        \cache_data_B[3][62] ) );
  dp_1 \cache_data_B_reg[3][63]  ( .ip(n5913), .ck(clk), .q(
        \cache_data_B[3][63] ) );
  dp_1 \cache_data_B_reg[4][32]  ( .ip(n5816), .ck(clk), .q(
        \cache_data_B[4][32] ) );
  dp_1 \cache_data_B_reg[4][33]  ( .ip(n5815), .ck(clk), .q(
        \cache_data_B[4][33] ) );
  dp_1 \cache_data_B_reg[4][34]  ( .ip(n5814), .ck(clk), .q(
        \cache_data_B[4][34] ) );
  dp_1 \cache_data_B_reg[4][35]  ( .ip(n5813), .ck(clk), .q(
        \cache_data_B[4][35] ) );
  dp_1 \cache_data_B_reg[4][36]  ( .ip(n5812), .ck(clk), .q(
        \cache_data_B[4][36] ) );
  dp_1 \cache_data_B_reg[4][37]  ( .ip(n5811), .ck(clk), .q(
        \cache_data_B[4][37] ) );
  dp_1 \cache_data_B_reg[4][38]  ( .ip(n5810), .ck(clk), .q(
        \cache_data_B[4][38] ) );
  dp_1 \cache_data_B_reg[4][39]  ( .ip(n5809), .ck(clk), .q(
        \cache_data_B[4][39] ) );
  dp_1 \cache_data_B_reg[4][40]  ( .ip(n5808), .ck(clk), .q(
        \cache_data_B[4][40] ) );
  dp_1 \cache_data_B_reg[4][41]  ( .ip(n5807), .ck(clk), .q(
        \cache_data_B[4][41] ) );
  dp_1 \cache_data_B_reg[4][42]  ( .ip(n5806), .ck(clk), .q(
        \cache_data_B[4][42] ) );
  dp_1 \cache_data_B_reg[4][43]  ( .ip(n5805), .ck(clk), .q(
        \cache_data_B[4][43] ) );
  dp_1 \cache_data_B_reg[4][44]  ( .ip(n5804), .ck(clk), .q(
        \cache_data_B[4][44] ) );
  dp_1 \cache_data_B_reg[4][45]  ( .ip(n5803), .ck(clk), .q(
        \cache_data_B[4][45] ) );
  dp_1 \cache_data_B_reg[4][46]  ( .ip(n5802), .ck(clk), .q(
        \cache_data_B[4][46] ) );
  dp_1 \cache_data_B_reg[4][47]  ( .ip(n5801), .ck(clk), .q(
        \cache_data_B[4][47] ) );
  dp_1 \cache_data_B_reg[4][48]  ( .ip(n5800), .ck(clk), .q(
        \cache_data_B[4][48] ) );
  dp_1 \cache_data_B_reg[4][49]  ( .ip(n5799), .ck(clk), .q(
        \cache_data_B[4][49] ) );
  dp_1 \cache_data_B_reg[4][50]  ( .ip(n5798), .ck(clk), .q(
        \cache_data_B[4][50] ) );
  dp_1 \cache_data_B_reg[4][51]  ( .ip(n5797), .ck(clk), .q(
        \cache_data_B[4][51] ) );
  dp_1 \cache_data_B_reg[4][52]  ( .ip(n5796), .ck(clk), .q(
        \cache_data_B[4][52] ) );
  dp_1 \cache_data_B_reg[4][53]  ( .ip(n5795), .ck(clk), .q(
        \cache_data_B[4][53] ) );
  dp_1 \cache_data_B_reg[4][54]  ( .ip(n5794), .ck(clk), .q(
        \cache_data_B[4][54] ) );
  dp_1 \cache_data_B_reg[4][55]  ( .ip(n5793), .ck(clk), .q(
        \cache_data_B[4][55] ) );
  dp_1 \cache_data_B_reg[4][56]  ( .ip(n5792), .ck(clk), .q(
        \cache_data_B[4][56] ) );
  dp_1 \cache_data_B_reg[4][57]  ( .ip(n5791), .ck(clk), .q(
        \cache_data_B[4][57] ) );
  dp_1 \cache_data_B_reg[4][58]  ( .ip(n5790), .ck(clk), .q(
        \cache_data_B[4][58] ) );
  dp_1 \cache_data_B_reg[4][59]  ( .ip(n5789), .ck(clk), .q(
        \cache_data_B[4][59] ) );
  dp_1 \cache_data_B_reg[4][60]  ( .ip(n5788), .ck(clk), .q(
        \cache_data_B[4][60] ) );
  dp_1 \cache_data_B_reg[4][61]  ( .ip(n5787), .ck(clk), .q(
        \cache_data_B[4][61] ) );
  dp_1 \cache_data_B_reg[4][62]  ( .ip(n5786), .ck(clk), .q(
        \cache_data_B[4][62] ) );
  dp_1 \cache_data_B_reg[4][63]  ( .ip(n5785), .ck(clk), .q(
        \cache_data_B[4][63] ) );
  dp_1 \cache_data_B_reg[5][42]  ( .ip(n5688), .ck(clk), .q(
        \cache_data_B[5][42] ) );
  dp_1 \cache_data_B_reg[5][43]  ( .ip(n5687), .ck(clk), .q(
        \cache_data_B[5][43] ) );
  dp_1 \cache_data_B_reg[5][44]  ( .ip(n5686), .ck(clk), .q(
        \cache_data_B[5][44] ) );
  dp_1 \cache_data_B_reg[5][45]  ( .ip(n5685), .ck(clk), .q(
        \cache_data_B[5][45] ) );
  dp_1 \cache_data_B_reg[5][46]  ( .ip(n5684), .ck(clk), .q(
        \cache_data_B[5][46] ) );
  dp_1 \cache_data_B_reg[5][47]  ( .ip(n5683), .ck(clk), .q(
        \cache_data_B[5][47] ) );
  dp_1 \cache_data_B_reg[5][48]  ( .ip(n5682), .ck(clk), .q(
        \cache_data_B[5][48] ) );
  dp_1 \cache_data_B_reg[5][49]  ( .ip(n5681), .ck(clk), .q(
        \cache_data_B[5][49] ) );
  dp_1 \cache_data_B_reg[5][50]  ( .ip(n5680), .ck(clk), .q(
        \cache_data_B[5][50] ) );
  dp_1 \cache_data_B_reg[5][51]  ( .ip(n5679), .ck(clk), .q(
        \cache_data_B[5][51] ) );
  dp_1 \cache_data_B_reg[5][52]  ( .ip(n5678), .ck(clk), .q(
        \cache_data_B[5][52] ) );
  dp_1 \cache_data_B_reg[5][53]  ( .ip(n5677), .ck(clk), .q(
        \cache_data_B[5][53] ) );
  dp_1 \cache_data_B_reg[5][54]  ( .ip(n5676), .ck(clk), .q(
        \cache_data_B[5][54] ) );
  dp_1 \cache_data_B_reg[5][55]  ( .ip(n5675), .ck(clk), .q(
        \cache_data_B[5][55] ) );
  dp_1 \cache_data_B_reg[5][56]  ( .ip(n5674), .ck(clk), .q(
        \cache_data_B[5][56] ) );
  dp_1 \cache_data_B_reg[5][57]  ( .ip(n5673), .ck(clk), .q(
        \cache_data_B[5][57] ) );
  dp_1 \cache_data_B_reg[5][58]  ( .ip(n5672), .ck(clk), .q(
        \cache_data_B[5][58] ) );
  dp_1 \cache_data_B_reg[5][59]  ( .ip(n5671), .ck(clk), .q(
        \cache_data_B[5][59] ) );
  dp_1 \cache_data_B_reg[5][60]  ( .ip(n5670), .ck(clk), .q(
        \cache_data_B[5][60] ) );
  dp_1 \cache_data_B_reg[5][61]  ( .ip(n5669), .ck(clk), .q(
        \cache_data_B[5][61] ) );
  dp_1 \cache_data_B_reg[5][62]  ( .ip(n5668), .ck(clk), .q(
        \cache_data_B[5][62] ) );
  dp_1 \cache_data_B_reg[5][63]  ( .ip(n5667), .ck(clk), .q(
        \cache_data_B[5][63] ) );
  dp_1 \cache_data_B_reg[5][32]  ( .ip(n5666), .ck(clk), .q(
        \cache_data_B[5][32] ) );
  dp_1 \cache_data_B_reg[5][33]  ( .ip(n5665), .ck(clk), .q(
        \cache_data_B[5][33] ) );
  dp_1 \cache_data_B_reg[5][34]  ( .ip(n5664), .ck(clk), .q(
        \cache_data_B[5][34] ) );
  dp_1 \cache_data_B_reg[5][35]  ( .ip(n5663), .ck(clk), .q(
        \cache_data_B[5][35] ) );
  dp_1 \cache_data_B_reg[5][36]  ( .ip(n5662), .ck(clk), .q(
        \cache_data_B[5][36] ) );
  dp_1 \cache_data_B_reg[5][37]  ( .ip(n5661), .ck(clk), .q(
        \cache_data_B[5][37] ) );
  dp_1 \cache_data_B_reg[5][38]  ( .ip(n5660), .ck(clk), .q(
        \cache_data_B[5][38] ) );
  dp_1 \cache_data_B_reg[5][39]  ( .ip(n5659), .ck(clk), .q(
        \cache_data_B[5][39] ) );
  dp_1 \cache_data_B_reg[5][40]  ( .ip(n5658), .ck(clk), .q(
        \cache_data_B[5][40] ) );
  dp_1 \cache_data_B_reg[5][41]  ( .ip(n5657), .ck(clk), .q(
        \cache_data_B[5][41] ) );
  dp_1 \cache_data_B_reg[6][32]  ( .ip(n5560), .ck(clk), .q(
        \cache_data_B[6][32] ) );
  dp_1 \cache_data_B_reg[6][33]  ( .ip(n5559), .ck(clk), .q(
        \cache_data_B[6][33] ) );
  dp_1 \cache_data_B_reg[6][34]  ( .ip(n5558), .ck(clk), .q(
        \cache_data_B[6][34] ) );
  dp_1 \cache_data_B_reg[6][35]  ( .ip(n5557), .ck(clk), .q(
        \cache_data_B[6][35] ) );
  dp_1 \cache_data_B_reg[6][36]  ( .ip(n5556), .ck(clk), .q(
        \cache_data_B[6][36] ) );
  dp_1 \cache_data_B_reg[6][37]  ( .ip(n5555), .ck(clk), .q(
        \cache_data_B[6][37] ) );
  dp_1 \cache_data_B_reg[6][38]  ( .ip(n5554), .ck(clk), .q(
        \cache_data_B[6][38] ) );
  dp_1 \cache_data_B_reg[6][39]  ( .ip(n5553), .ck(clk), .q(
        \cache_data_B[6][39] ) );
  dp_1 \cache_data_B_reg[6][40]  ( .ip(n5552), .ck(clk), .q(
        \cache_data_B[6][40] ) );
  dp_1 \cache_data_B_reg[6][41]  ( .ip(n5551), .ck(clk), .q(
        \cache_data_B[6][41] ) );
  dp_1 \cache_data_B_reg[6][42]  ( .ip(n5550), .ck(clk), .q(
        \cache_data_B[6][42] ) );
  dp_1 \cache_data_B_reg[6][43]  ( .ip(n5549), .ck(clk), .q(
        \cache_data_B[6][43] ) );
  dp_1 \cache_data_B_reg[6][44]  ( .ip(n5548), .ck(clk), .q(
        \cache_data_B[6][44] ) );
  dp_1 \cache_data_B_reg[6][45]  ( .ip(n5547), .ck(clk), .q(
        \cache_data_B[6][45] ) );
  dp_1 \cache_data_B_reg[6][46]  ( .ip(n5546), .ck(clk), .q(
        \cache_data_B[6][46] ) );
  dp_1 \cache_data_B_reg[6][47]  ( .ip(n5545), .ck(clk), .q(
        \cache_data_B[6][47] ) );
  dp_1 \cache_data_B_reg[6][48]  ( .ip(n5544), .ck(clk), .q(
        \cache_data_B[6][48] ) );
  dp_1 \cache_data_B_reg[6][49]  ( .ip(n5543), .ck(clk), .q(
        \cache_data_B[6][49] ) );
  dp_1 \cache_data_B_reg[6][50]  ( .ip(n5542), .ck(clk), .q(
        \cache_data_B[6][50] ) );
  dp_1 \cache_data_B_reg[6][51]  ( .ip(n5541), .ck(clk), .q(
        \cache_data_B[6][51] ) );
  dp_1 \cache_data_B_reg[6][52]  ( .ip(n5540), .ck(clk), .q(
        \cache_data_B[6][52] ) );
  dp_1 \cache_data_B_reg[6][53]  ( .ip(n5539), .ck(clk), .q(
        \cache_data_B[6][53] ) );
  dp_1 \cache_data_B_reg[6][54]  ( .ip(n5538), .ck(clk), .q(
        \cache_data_B[6][54] ) );
  dp_1 \cache_data_B_reg[6][55]  ( .ip(n5537), .ck(clk), .q(
        \cache_data_B[6][55] ) );
  dp_1 \cache_data_B_reg[6][56]  ( .ip(n5536), .ck(clk), .q(
        \cache_data_B[6][56] ) );
  dp_1 \cache_data_B_reg[6][57]  ( .ip(n5535), .ck(clk), .q(
        \cache_data_B[6][57] ) );
  dp_1 \cache_data_B_reg[6][58]  ( .ip(n5534), .ck(clk), .q(
        \cache_data_B[6][58] ) );
  dp_1 \cache_data_B_reg[6][59]  ( .ip(n5533), .ck(clk), .q(
        \cache_data_B[6][59] ) );
  dp_1 \cache_data_B_reg[6][60]  ( .ip(n5532), .ck(clk), .q(
        \cache_data_B[6][60] ) );
  dp_1 \cache_data_B_reg[6][61]  ( .ip(n5531), .ck(clk), .q(
        \cache_data_B[6][61] ) );
  dp_1 \cache_data_B_reg[6][62]  ( .ip(n5530), .ck(clk), .q(
        \cache_data_B[6][62] ) );
  dp_1 \cache_data_B_reg[6][63]  ( .ip(n5529), .ck(clk), .q(
        \cache_data_B[6][63] ) );
  dp_1 \cache_data_B_reg[7][32]  ( .ip(n5432), .ck(clk), .q(
        \cache_data_B[7][32] ) );
  dp_1 \cache_data_B_reg[7][33]  ( .ip(n5431), .ck(clk), .q(
        \cache_data_B[7][33] ) );
  dp_1 \cache_data_B_reg[7][34]  ( .ip(n5430), .ck(clk), .q(
        \cache_data_B[7][34] ) );
  dp_1 \cache_data_B_reg[7][35]  ( .ip(n5429), .ck(clk), .q(
        \cache_data_B[7][35] ) );
  dp_1 \cache_data_B_reg[7][36]  ( .ip(n5428), .ck(clk), .q(
        \cache_data_B[7][36] ) );
  dp_1 \cache_data_B_reg[7][37]  ( .ip(n5427), .ck(clk), .q(
        \cache_data_B[7][37] ) );
  dp_1 \cache_data_B_reg[7][38]  ( .ip(n5426), .ck(clk), .q(
        \cache_data_B[7][38] ) );
  dp_1 \cache_data_B_reg[7][39]  ( .ip(n5425), .ck(clk), .q(
        \cache_data_B[7][39] ) );
  dp_1 \cache_data_B_reg[7][40]  ( .ip(n5424), .ck(clk), .q(
        \cache_data_B[7][40] ) );
  dp_1 \cache_data_B_reg[7][41]  ( .ip(n5423), .ck(clk), .q(
        \cache_data_B[7][41] ) );
  dp_1 \cache_data_B_reg[7][42]  ( .ip(n5422), .ck(clk), .q(
        \cache_data_B[7][42] ) );
  dp_1 \cache_data_B_reg[7][43]  ( .ip(n5421), .ck(clk), .q(
        \cache_data_B[7][43] ) );
  dp_1 \cache_data_B_reg[7][44]  ( .ip(n5420), .ck(clk), .q(
        \cache_data_B[7][44] ) );
  dp_1 \cache_data_B_reg[7][45]  ( .ip(n5419), .ck(clk), .q(
        \cache_data_B[7][45] ) );
  dp_1 \cache_data_B_reg[7][46]  ( .ip(n5418), .ck(clk), .q(
        \cache_data_B[7][46] ) );
  dp_1 \cache_data_B_reg[7][47]  ( .ip(n5417), .ck(clk), .q(
        \cache_data_B[7][47] ) );
  dp_1 \cache_data_B_reg[7][48]  ( .ip(n5416), .ck(clk), .q(
        \cache_data_B[7][48] ) );
  dp_1 \cache_data_B_reg[7][49]  ( .ip(n5415), .ck(clk), .q(
        \cache_data_B[7][49] ) );
  dp_1 \cache_data_B_reg[7][50]  ( .ip(n5414), .ck(clk), .q(
        \cache_data_B[7][50] ) );
  dp_1 \cache_data_B_reg[7][51]  ( .ip(n5413), .ck(clk), .q(
        \cache_data_B[7][51] ) );
  dp_1 \cache_data_B_reg[7][52]  ( .ip(n5412), .ck(clk), .q(
        \cache_data_B[7][52] ) );
  dp_1 \cache_data_B_reg[7][53]  ( .ip(n5411), .ck(clk), .q(
        \cache_data_B[7][53] ) );
  dp_1 \cache_data_B_reg[7][54]  ( .ip(n5410), .ck(clk), .q(
        \cache_data_B[7][54] ) );
  dp_1 \cache_data_B_reg[7][55]  ( .ip(n5409), .ck(clk), .q(
        \cache_data_B[7][55] ) );
  dp_1 \cache_data_B_reg[7][56]  ( .ip(n5408), .ck(clk), .q(
        \cache_data_B[7][56] ) );
  dp_1 \cache_data_B_reg[7][57]  ( .ip(n5407), .ck(clk), .q(
        \cache_data_B[7][57] ) );
  dp_1 \cache_data_B_reg[7][58]  ( .ip(n5406), .ck(clk), .q(
        \cache_data_B[7][58] ) );
  dp_1 \cache_data_B_reg[7][59]  ( .ip(n5405), .ck(clk), .q(
        \cache_data_B[7][59] ) );
  dp_1 \cache_data_B_reg[7][60]  ( .ip(n5404), .ck(clk), .q(
        \cache_data_B[7][60] ) );
  dp_1 \cache_data_B_reg[7][61]  ( .ip(n5403), .ck(clk), .q(
        \cache_data_B[7][61] ) );
  dp_1 \cache_data_B_reg[7][62]  ( .ip(n5402), .ck(clk), .q(
        \cache_data_B[7][62] ) );
  dp_1 \cache_data_B_reg[7][63]  ( .ip(n5401), .ck(clk), .q(
        \cache_data_B[7][63] ) );
  dp_1 \cache_data_B_reg[0][88]  ( .ip(n6296), .ck(clk), .q(
        \cache_data_B[0][88] ) );
  dp_1 \cache_data_B_reg[0][89]  ( .ip(n6295), .ck(clk), .q(
        \cache_data_B[0][89] ) );
  dp_1 \cache_data_B_reg[0][90]  ( .ip(n6294), .ck(clk), .q(
        \cache_data_B[0][90] ) );
  dp_1 \cache_data_B_reg[0][91]  ( .ip(n6293), .ck(clk), .q(
        \cache_data_B[0][91] ) );
  dp_1 \cache_data_B_reg[0][92]  ( .ip(n6292), .ck(clk), .q(
        \cache_data_B[0][92] ) );
  dp_1 \cache_data_B_reg[0][93]  ( .ip(n6291), .ck(clk), .q(
        \cache_data_B[0][93] ) );
  dp_1 \cache_data_B_reg[0][94]  ( .ip(n6290), .ck(clk), .q(
        \cache_data_B[0][94] ) );
  dp_1 \cache_data_B_reg[0][95]  ( .ip(n6289), .ck(clk), .q(
        \cache_data_B[0][95] ) );
  dp_1 \cache_data_B_reg[0][64]  ( .ip(n6288), .ck(clk), .q(
        \cache_data_B[0][64] ) );
  dp_1 \cache_data_B_reg[0][65]  ( .ip(n6287), .ck(clk), .q(
        \cache_data_B[0][65] ) );
  dp_1 \cache_data_B_reg[0][66]  ( .ip(n6286), .ck(clk), .q(
        \cache_data_B[0][66] ) );
  dp_1 \cache_data_B_reg[0][67]  ( .ip(n6285), .ck(clk), .q(
        \cache_data_B[0][67] ) );
  dp_1 \cache_data_B_reg[0][68]  ( .ip(n6284), .ck(clk), .q(
        \cache_data_B[0][68] ) );
  dp_1 \cache_data_B_reg[0][69]  ( .ip(n6283), .ck(clk), .q(
        \cache_data_B[0][69] ) );
  dp_1 \cache_data_B_reg[0][70]  ( .ip(n6282), .ck(clk), .q(
        \cache_data_B[0][70] ) );
  dp_1 \cache_data_B_reg[0][71]  ( .ip(n6281), .ck(clk), .q(
        \cache_data_B[0][71] ) );
  dp_1 \cache_data_B_reg[0][72]  ( .ip(n6280), .ck(clk), .q(
        \cache_data_B[0][72] ) );
  dp_1 \cache_data_B_reg[0][73]  ( .ip(n6279), .ck(clk), .q(
        \cache_data_B[0][73] ) );
  dp_1 \cache_data_B_reg[0][74]  ( .ip(n6278), .ck(clk), .q(
        \cache_data_B[0][74] ) );
  dp_1 \cache_data_B_reg[0][75]  ( .ip(n6277), .ck(clk), .q(
        \cache_data_B[0][75] ) );
  dp_1 \cache_data_B_reg[0][76]  ( .ip(n6276), .ck(clk), .q(
        \cache_data_B[0][76] ) );
  dp_1 \cache_data_B_reg[0][77]  ( .ip(n6275), .ck(clk), .q(
        \cache_data_B[0][77] ) );
  dp_1 \cache_data_B_reg[0][78]  ( .ip(n6274), .ck(clk), .q(
        \cache_data_B[0][78] ) );
  dp_1 \cache_data_B_reg[0][79]  ( .ip(n6273), .ck(clk), .q(
        \cache_data_B[0][79] ) );
  dp_1 \cache_data_B_reg[0][80]  ( .ip(n6272), .ck(clk), .q(
        \cache_data_B[0][80] ) );
  dp_1 \cache_data_B_reg[0][81]  ( .ip(n6271), .ck(clk), .q(
        \cache_data_B[0][81] ) );
  dp_1 \cache_data_B_reg[0][82]  ( .ip(n6270), .ck(clk), .q(
        \cache_data_B[0][82] ) );
  dp_1 \cache_data_B_reg[0][83]  ( .ip(n6269), .ck(clk), .q(
        \cache_data_B[0][83] ) );
  dp_1 \cache_data_B_reg[0][84]  ( .ip(n6268), .ck(clk), .q(
        \cache_data_B[0][84] ) );
  dp_1 \cache_data_B_reg[0][85]  ( .ip(n6267), .ck(clk), .q(
        \cache_data_B[0][85] ) );
  dp_1 \cache_data_B_reg[0][86]  ( .ip(n6266), .ck(clk), .q(
        \cache_data_B[0][86] ) );
  dp_1 \cache_data_B_reg[0][87]  ( .ip(n6265), .ck(clk), .q(
        \cache_data_B[0][87] ) );
  dp_1 \cache_data_B_reg[1][64]  ( .ip(n6168), .ck(clk), .q(
        \cache_data_B[1][64] ) );
  dp_1 \cache_data_B_reg[1][65]  ( .ip(n6167), .ck(clk), .q(
        \cache_data_B[1][65] ) );
  dp_1 \cache_data_B_reg[1][66]  ( .ip(n6166), .ck(clk), .q(
        \cache_data_B[1][66] ) );
  dp_1 \cache_data_B_reg[1][67]  ( .ip(n6165), .ck(clk), .q(
        \cache_data_B[1][67] ) );
  dp_1 \cache_data_B_reg[1][68]  ( .ip(n6164), .ck(clk), .q(
        \cache_data_B[1][68] ) );
  dp_1 \cache_data_B_reg[1][69]  ( .ip(n6163), .ck(clk), .q(
        \cache_data_B[1][69] ) );
  dp_1 \cache_data_B_reg[1][70]  ( .ip(n6162), .ck(clk), .q(
        \cache_data_B[1][70] ) );
  dp_1 \cache_data_B_reg[1][71]  ( .ip(n6161), .ck(clk), .q(
        \cache_data_B[1][71] ) );
  dp_1 \cache_data_B_reg[1][72]  ( .ip(n6160), .ck(clk), .q(
        \cache_data_B[1][72] ) );
  dp_1 \cache_data_B_reg[1][73]  ( .ip(n6159), .ck(clk), .q(
        \cache_data_B[1][73] ) );
  dp_1 \cache_data_B_reg[1][74]  ( .ip(n6158), .ck(clk), .q(
        \cache_data_B[1][74] ) );
  dp_1 \cache_data_B_reg[1][75]  ( .ip(n6157), .ck(clk), .q(
        \cache_data_B[1][75] ) );
  dp_1 \cache_data_B_reg[1][76]  ( .ip(n6156), .ck(clk), .q(
        \cache_data_B[1][76] ) );
  dp_1 \cache_data_B_reg[1][77]  ( .ip(n6155), .ck(clk), .q(
        \cache_data_B[1][77] ) );
  dp_1 \cache_data_B_reg[1][78]  ( .ip(n6154), .ck(clk), .q(
        \cache_data_B[1][78] ) );
  dp_1 \cache_data_B_reg[1][79]  ( .ip(n6153), .ck(clk), .q(
        \cache_data_B[1][79] ) );
  dp_1 \cache_data_B_reg[1][80]  ( .ip(n6152), .ck(clk), .q(
        \cache_data_B[1][80] ) );
  dp_1 \cache_data_B_reg[1][81]  ( .ip(n6151), .ck(clk), .q(
        \cache_data_B[1][81] ) );
  dp_1 \cache_data_B_reg[1][82]  ( .ip(n6150), .ck(clk), .q(
        \cache_data_B[1][82] ) );
  dp_1 \cache_data_B_reg[1][83]  ( .ip(n6149), .ck(clk), .q(
        \cache_data_B[1][83] ) );
  dp_1 \cache_data_B_reg[1][84]  ( .ip(n6148), .ck(clk), .q(
        \cache_data_B[1][84] ) );
  dp_1 \cache_data_B_reg[1][85]  ( .ip(n6147), .ck(clk), .q(
        \cache_data_B[1][85] ) );
  dp_1 \cache_data_B_reg[1][86]  ( .ip(n6146), .ck(clk), .q(
        \cache_data_B[1][86] ) );
  dp_1 \cache_data_B_reg[1][87]  ( .ip(n6145), .ck(clk), .q(
        \cache_data_B[1][87] ) );
  dp_1 \cache_data_B_reg[1][88]  ( .ip(n6144), .ck(clk), .q(
        \cache_data_B[1][88] ) );
  dp_1 \cache_data_B_reg[1][89]  ( .ip(n6143), .ck(clk), .q(
        \cache_data_B[1][89] ) );
  dp_1 \cache_data_B_reg[1][90]  ( .ip(n6142), .ck(clk), .q(
        \cache_data_B[1][90] ) );
  dp_1 \cache_data_B_reg[1][91]  ( .ip(n6141), .ck(clk), .q(
        \cache_data_B[1][91] ) );
  dp_1 \cache_data_B_reg[1][92]  ( .ip(n6140), .ck(clk), .q(
        \cache_data_B[1][92] ) );
  dp_1 \cache_data_B_reg[1][93]  ( .ip(n6139), .ck(clk), .q(
        \cache_data_B[1][93] ) );
  dp_1 \cache_data_B_reg[1][94]  ( .ip(n6138), .ck(clk), .q(
        \cache_data_B[1][94] ) );
  dp_1 \cache_data_B_reg[1][95]  ( .ip(n6137), .ck(clk), .q(
        \cache_data_B[1][95] ) );
  dp_1 \cache_data_B_reg[2][64]  ( .ip(n6040), .ck(clk), .q(
        \cache_data_B[2][64] ) );
  dp_1 \cache_data_B_reg[2][65]  ( .ip(n6039), .ck(clk), .q(
        \cache_data_B[2][65] ) );
  dp_1 \cache_data_B_reg[2][66]  ( .ip(n6038), .ck(clk), .q(
        \cache_data_B[2][66] ) );
  dp_1 \cache_data_B_reg[2][67]  ( .ip(n6037), .ck(clk), .q(
        \cache_data_B[2][67] ) );
  dp_1 \cache_data_B_reg[2][68]  ( .ip(n6036), .ck(clk), .q(
        \cache_data_B[2][68] ) );
  dp_1 \cache_data_B_reg[2][69]  ( .ip(n6035), .ck(clk), .q(
        \cache_data_B[2][69] ) );
  dp_1 \cache_data_B_reg[2][70]  ( .ip(n6034), .ck(clk), .q(
        \cache_data_B[2][70] ) );
  dp_1 \cache_data_B_reg[2][71]  ( .ip(n6033), .ck(clk), .q(
        \cache_data_B[2][71] ) );
  dp_1 \cache_data_B_reg[2][72]  ( .ip(n6032), .ck(clk), .q(
        \cache_data_B[2][72] ) );
  dp_1 \cache_data_B_reg[2][73]  ( .ip(n6031), .ck(clk), .q(
        \cache_data_B[2][73] ) );
  dp_1 \cache_data_B_reg[2][74]  ( .ip(n6030), .ck(clk), .q(
        \cache_data_B[2][74] ) );
  dp_1 \cache_data_B_reg[2][75]  ( .ip(n6029), .ck(clk), .q(
        \cache_data_B[2][75] ) );
  dp_1 \cache_data_B_reg[2][76]  ( .ip(n6028), .ck(clk), .q(
        \cache_data_B[2][76] ) );
  dp_1 \cache_data_B_reg[2][77]  ( .ip(n6027), .ck(clk), .q(
        \cache_data_B[2][77] ) );
  dp_1 \cache_data_B_reg[2][78]  ( .ip(n6026), .ck(clk), .q(
        \cache_data_B[2][78] ) );
  dp_1 \cache_data_B_reg[2][79]  ( .ip(n6025), .ck(clk), .q(
        \cache_data_B[2][79] ) );
  dp_1 \cache_data_B_reg[2][80]  ( .ip(n6024), .ck(clk), .q(
        \cache_data_B[2][80] ) );
  dp_1 \cache_data_B_reg[2][81]  ( .ip(n6023), .ck(clk), .q(
        \cache_data_B[2][81] ) );
  dp_1 \cache_data_B_reg[2][82]  ( .ip(n6022), .ck(clk), .q(
        \cache_data_B[2][82] ) );
  dp_1 \cache_data_B_reg[2][83]  ( .ip(n6021), .ck(clk), .q(
        \cache_data_B[2][83] ) );
  dp_1 \cache_data_B_reg[2][84]  ( .ip(n6020), .ck(clk), .q(
        \cache_data_B[2][84] ) );
  dp_1 \cache_data_B_reg[2][85]  ( .ip(n6019), .ck(clk), .q(
        \cache_data_B[2][85] ) );
  dp_1 \cache_data_B_reg[2][86]  ( .ip(n6018), .ck(clk), .q(
        \cache_data_B[2][86] ) );
  dp_1 \cache_data_B_reg[2][87]  ( .ip(n6017), .ck(clk), .q(
        \cache_data_B[2][87] ) );
  dp_1 \cache_data_B_reg[2][88]  ( .ip(n6016), .ck(clk), .q(
        \cache_data_B[2][88] ) );
  dp_1 \cache_data_B_reg[2][89]  ( .ip(n6015), .ck(clk), .q(
        \cache_data_B[2][89] ) );
  dp_1 \cache_data_B_reg[2][90]  ( .ip(n6014), .ck(clk), .q(
        \cache_data_B[2][90] ) );
  dp_1 \cache_data_B_reg[2][91]  ( .ip(n6013), .ck(clk), .q(
        \cache_data_B[2][91] ) );
  dp_1 \cache_data_B_reg[2][92]  ( .ip(n6012), .ck(clk), .q(
        \cache_data_B[2][92] ) );
  dp_1 \cache_data_B_reg[2][93]  ( .ip(n6011), .ck(clk), .q(
        \cache_data_B[2][93] ) );
  dp_1 \cache_data_B_reg[2][94]  ( .ip(n6010), .ck(clk), .q(
        \cache_data_B[2][94] ) );
  dp_1 \cache_data_B_reg[2][95]  ( .ip(n6009), .ck(clk), .q(
        \cache_data_B[2][95] ) );
  dp_1 \cache_data_B_reg[3][64]  ( .ip(n5912), .ck(clk), .q(
        \cache_data_B[3][64] ) );
  dp_1 \cache_data_B_reg[3][65]  ( .ip(n5911), .ck(clk), .q(
        \cache_data_B[3][65] ) );
  dp_1 \cache_data_B_reg[3][66]  ( .ip(n5910), .ck(clk), .q(
        \cache_data_B[3][66] ) );
  dp_1 \cache_data_B_reg[3][67]  ( .ip(n5909), .ck(clk), .q(
        \cache_data_B[3][67] ) );
  dp_1 \cache_data_B_reg[3][68]  ( .ip(n5908), .ck(clk), .q(
        \cache_data_B[3][68] ) );
  dp_1 \cache_data_B_reg[3][69]  ( .ip(n5907), .ck(clk), .q(
        \cache_data_B[3][69] ) );
  dp_1 \cache_data_B_reg[3][70]  ( .ip(n5906), .ck(clk), .q(
        \cache_data_B[3][70] ) );
  dp_1 \cache_data_B_reg[3][71]  ( .ip(n5905), .ck(clk), .q(
        \cache_data_B[3][71] ) );
  dp_1 \cache_data_B_reg[3][72]  ( .ip(n5904), .ck(clk), .q(
        \cache_data_B[3][72] ) );
  dp_1 \cache_data_B_reg[3][73]  ( .ip(n5903), .ck(clk), .q(
        \cache_data_B[3][73] ) );
  dp_1 \cache_data_B_reg[3][74]  ( .ip(n5902), .ck(clk), .q(
        \cache_data_B[3][74] ) );
  dp_1 \cache_data_B_reg[3][75]  ( .ip(n5901), .ck(clk), .q(
        \cache_data_B[3][75] ) );
  dp_1 \cache_data_B_reg[3][76]  ( .ip(n5900), .ck(clk), .q(
        \cache_data_B[3][76] ) );
  dp_1 \cache_data_B_reg[3][77]  ( .ip(n5899), .ck(clk), .q(
        \cache_data_B[3][77] ) );
  dp_1 \cache_data_B_reg[3][78]  ( .ip(n5898), .ck(clk), .q(
        \cache_data_B[3][78] ) );
  dp_1 \cache_data_B_reg[3][79]  ( .ip(n5897), .ck(clk), .q(
        \cache_data_B[3][79] ) );
  dp_1 \cache_data_B_reg[3][80]  ( .ip(n5896), .ck(clk), .q(
        \cache_data_B[3][80] ) );
  dp_1 \cache_data_B_reg[3][81]  ( .ip(n5895), .ck(clk), .q(
        \cache_data_B[3][81] ) );
  dp_1 \cache_data_B_reg[3][82]  ( .ip(n5894), .ck(clk), .q(
        \cache_data_B[3][82] ) );
  dp_1 \cache_data_B_reg[3][83]  ( .ip(n5893), .ck(clk), .q(
        \cache_data_B[3][83] ) );
  dp_1 \cache_data_B_reg[3][84]  ( .ip(n5892), .ck(clk), .q(
        \cache_data_B[3][84] ) );
  dp_1 \cache_data_B_reg[3][85]  ( .ip(n5891), .ck(clk), .q(
        \cache_data_B[3][85] ) );
  dp_1 \cache_data_B_reg[3][86]  ( .ip(n5890), .ck(clk), .q(
        \cache_data_B[3][86] ) );
  dp_1 \cache_data_B_reg[3][87]  ( .ip(n5889), .ck(clk), .q(
        \cache_data_B[3][87] ) );
  dp_1 \cache_data_B_reg[3][88]  ( .ip(n5888), .ck(clk), .q(
        \cache_data_B[3][88] ) );
  dp_1 \cache_data_B_reg[3][89]  ( .ip(n5887), .ck(clk), .q(
        \cache_data_B[3][89] ) );
  dp_1 \cache_data_B_reg[3][90]  ( .ip(n5886), .ck(clk), .q(
        \cache_data_B[3][90] ) );
  dp_1 \cache_data_B_reg[3][91]  ( .ip(n5885), .ck(clk), .q(
        \cache_data_B[3][91] ) );
  dp_1 \cache_data_B_reg[3][92]  ( .ip(n5884), .ck(clk), .q(
        \cache_data_B[3][92] ) );
  dp_1 \cache_data_B_reg[3][93]  ( .ip(n5883), .ck(clk), .q(
        \cache_data_B[3][93] ) );
  dp_1 \cache_data_B_reg[3][94]  ( .ip(n5882), .ck(clk), .q(
        \cache_data_B[3][94] ) );
  dp_1 \cache_data_B_reg[3][95]  ( .ip(n5881), .ck(clk), .q(
        \cache_data_B[3][95] ) );
  dp_1 \cache_data_B_reg[4][71]  ( .ip(n5784), .ck(clk), .q(
        \cache_data_B[4][71] ) );
  dp_1 \cache_data_B_reg[4][72]  ( .ip(n5783), .ck(clk), .q(
        \cache_data_B[4][72] ) );
  dp_1 \cache_data_B_reg[4][73]  ( .ip(n5782), .ck(clk), .q(
        \cache_data_B[4][73] ) );
  dp_1 \cache_data_B_reg[4][74]  ( .ip(n5781), .ck(clk), .q(
        \cache_data_B[4][74] ) );
  dp_1 \cache_data_B_reg[4][75]  ( .ip(n5780), .ck(clk), .q(
        \cache_data_B[4][75] ) );
  dp_1 \cache_data_B_reg[4][76]  ( .ip(n5779), .ck(clk), .q(
        \cache_data_B[4][76] ) );
  dp_1 \cache_data_B_reg[4][77]  ( .ip(n5778), .ck(clk), .q(
        \cache_data_B[4][77] ) );
  dp_1 \cache_data_B_reg[4][78]  ( .ip(n5777), .ck(clk), .q(
        \cache_data_B[4][78] ) );
  dp_1 \cache_data_B_reg[4][79]  ( .ip(n5776), .ck(clk), .q(
        \cache_data_B[4][79] ) );
  dp_1 \cache_data_B_reg[4][80]  ( .ip(n5775), .ck(clk), .q(
        \cache_data_B[4][80] ) );
  dp_1 \cache_data_B_reg[4][81]  ( .ip(n5774), .ck(clk), .q(
        \cache_data_B[4][81] ) );
  dp_1 \cache_data_B_reg[4][82]  ( .ip(n5773), .ck(clk), .q(
        \cache_data_B[4][82] ) );
  dp_1 \cache_data_B_reg[4][83]  ( .ip(n5772), .ck(clk), .q(
        \cache_data_B[4][83] ) );
  dp_1 \cache_data_B_reg[4][84]  ( .ip(n5771), .ck(clk), .q(
        \cache_data_B[4][84] ) );
  dp_1 \cache_data_B_reg[4][85]  ( .ip(n5770), .ck(clk), .q(
        \cache_data_B[4][85] ) );
  dp_1 \cache_data_B_reg[4][86]  ( .ip(n5769), .ck(clk), .q(
        \cache_data_B[4][86] ) );
  dp_1 \cache_data_B_reg[4][87]  ( .ip(n5768), .ck(clk), .q(
        \cache_data_B[4][87] ) );
  dp_1 \cache_data_B_reg[4][88]  ( .ip(n5767), .ck(clk), .q(
        \cache_data_B[4][88] ) );
  dp_1 \cache_data_B_reg[4][89]  ( .ip(n5766), .ck(clk), .q(
        \cache_data_B[4][89] ) );
  dp_1 \cache_data_B_reg[4][90]  ( .ip(n5765), .ck(clk), .q(
        \cache_data_B[4][90] ) );
  dp_1 \cache_data_B_reg[4][91]  ( .ip(n5764), .ck(clk), .q(
        \cache_data_B[4][91] ) );
  dp_1 \cache_data_B_reg[4][92]  ( .ip(n5763), .ck(clk), .q(
        \cache_data_B[4][92] ) );
  dp_1 \cache_data_B_reg[4][93]  ( .ip(n5762), .ck(clk), .q(
        \cache_data_B[4][93] ) );
  dp_1 \cache_data_B_reg[4][94]  ( .ip(n5761), .ck(clk), .q(
        \cache_data_B[4][94] ) );
  dp_1 \cache_data_B_reg[4][95]  ( .ip(n5760), .ck(clk), .q(
        \cache_data_B[4][95] ) );
  dp_1 \cache_data_B_reg[4][64]  ( .ip(n5759), .ck(clk), .q(
        \cache_data_B[4][64] ) );
  dp_1 \cache_data_B_reg[4][65]  ( .ip(n5758), .ck(clk), .q(
        \cache_data_B[4][65] ) );
  dp_1 \cache_data_B_reg[4][66]  ( .ip(n5757), .ck(clk), .q(
        \cache_data_B[4][66] ) );
  dp_1 \cache_data_B_reg[4][67]  ( .ip(n5756), .ck(clk), .q(
        \cache_data_B[4][67] ) );
  dp_1 \cache_data_B_reg[4][68]  ( .ip(n5755), .ck(clk), .q(
        \cache_data_B[4][68] ) );
  dp_1 \cache_data_B_reg[4][69]  ( .ip(n5754), .ck(clk), .q(
        \cache_data_B[4][69] ) );
  dp_1 \cache_data_B_reg[4][70]  ( .ip(n5753), .ck(clk), .q(
        \cache_data_B[4][70] ) );
  dp_1 \cache_data_B_reg[5][64]  ( .ip(n5656), .ck(clk), .q(
        \cache_data_B[5][64] ) );
  dp_1 \cache_data_B_reg[5][65]  ( .ip(n5655), .ck(clk), .q(
        \cache_data_B[5][65] ) );
  dp_1 \cache_data_B_reg[5][66]  ( .ip(n5654), .ck(clk), .q(
        \cache_data_B[5][66] ) );
  dp_1 \cache_data_B_reg[5][67]  ( .ip(n5653), .ck(clk), .q(
        \cache_data_B[5][67] ) );
  dp_1 \cache_data_B_reg[5][68]  ( .ip(n5652), .ck(clk), .q(
        \cache_data_B[5][68] ) );
  dp_1 \cache_data_B_reg[5][69]  ( .ip(n5651), .ck(clk), .q(
        \cache_data_B[5][69] ) );
  dp_1 \cache_data_B_reg[5][70]  ( .ip(n5650), .ck(clk), .q(
        \cache_data_B[5][70] ) );
  dp_1 \cache_data_B_reg[5][71]  ( .ip(n5649), .ck(clk), .q(
        \cache_data_B[5][71] ) );
  dp_1 \cache_data_B_reg[5][72]  ( .ip(n5648), .ck(clk), .q(
        \cache_data_B[5][72] ) );
  dp_1 \cache_data_B_reg[5][73]  ( .ip(n5647), .ck(clk), .q(
        \cache_data_B[5][73] ) );
  dp_1 \cache_data_B_reg[5][74]  ( .ip(n5646), .ck(clk), .q(
        \cache_data_B[5][74] ) );
  dp_1 \cache_data_B_reg[5][75]  ( .ip(n5645), .ck(clk), .q(
        \cache_data_B[5][75] ) );
  dp_1 \cache_data_B_reg[5][76]  ( .ip(n5644), .ck(clk), .q(
        \cache_data_B[5][76] ) );
  dp_1 \cache_data_B_reg[5][77]  ( .ip(n5643), .ck(clk), .q(
        \cache_data_B[5][77] ) );
  dp_1 \cache_data_B_reg[5][78]  ( .ip(n5642), .ck(clk), .q(
        \cache_data_B[5][78] ) );
  dp_1 \cache_data_B_reg[5][79]  ( .ip(n5641), .ck(clk), .q(
        \cache_data_B[5][79] ) );
  dp_1 \cache_data_B_reg[5][80]  ( .ip(n5640), .ck(clk), .q(
        \cache_data_B[5][80] ) );
  dp_1 \cache_data_B_reg[5][81]  ( .ip(n5639), .ck(clk), .q(
        \cache_data_B[5][81] ) );
  dp_1 \cache_data_B_reg[5][82]  ( .ip(n5638), .ck(clk), .q(
        \cache_data_B[5][82] ) );
  dp_1 \cache_data_B_reg[5][83]  ( .ip(n5637), .ck(clk), .q(
        \cache_data_B[5][83] ) );
  dp_1 \cache_data_B_reg[5][84]  ( .ip(n5636), .ck(clk), .q(
        \cache_data_B[5][84] ) );
  dp_1 \cache_data_B_reg[5][85]  ( .ip(n5635), .ck(clk), .q(
        \cache_data_B[5][85] ) );
  dp_1 \cache_data_B_reg[5][86]  ( .ip(n5634), .ck(clk), .q(
        \cache_data_B[5][86] ) );
  dp_1 \cache_data_B_reg[5][87]  ( .ip(n5633), .ck(clk), .q(
        \cache_data_B[5][87] ) );
  dp_1 \cache_data_B_reg[5][88]  ( .ip(n5632), .ck(clk), .q(
        \cache_data_B[5][88] ) );
  dp_1 \cache_data_B_reg[5][89]  ( .ip(n5631), .ck(clk), .q(
        \cache_data_B[5][89] ) );
  dp_1 \cache_data_B_reg[5][90]  ( .ip(n5630), .ck(clk), .q(
        \cache_data_B[5][90] ) );
  dp_1 \cache_data_B_reg[5][91]  ( .ip(n5629), .ck(clk), .q(
        \cache_data_B[5][91] ) );
  dp_1 \cache_data_B_reg[5][92]  ( .ip(n5628), .ck(clk), .q(
        \cache_data_B[5][92] ) );
  dp_1 \cache_data_B_reg[5][93]  ( .ip(n5627), .ck(clk), .q(
        \cache_data_B[5][93] ) );
  dp_1 \cache_data_B_reg[5][94]  ( .ip(n5626), .ck(clk), .q(
        \cache_data_B[5][94] ) );
  dp_1 \cache_data_B_reg[5][95]  ( .ip(n5625), .ck(clk), .q(
        \cache_data_B[5][95] ) );
  dp_1 \cache_data_B_reg[6][64]  ( .ip(n5528), .ck(clk), .q(
        \cache_data_B[6][64] ) );
  dp_1 \cache_data_B_reg[6][65]  ( .ip(n5527), .ck(clk), .q(
        \cache_data_B[6][65] ) );
  dp_1 \cache_data_B_reg[6][66]  ( .ip(n5526), .ck(clk), .q(
        \cache_data_B[6][66] ) );
  dp_1 \cache_data_B_reg[6][67]  ( .ip(n5525), .ck(clk), .q(
        \cache_data_B[6][67] ) );
  dp_1 \cache_data_B_reg[6][68]  ( .ip(n5524), .ck(clk), .q(
        \cache_data_B[6][68] ) );
  dp_1 \cache_data_B_reg[6][69]  ( .ip(n5523), .ck(clk), .q(
        \cache_data_B[6][69] ) );
  dp_1 \cache_data_B_reg[6][70]  ( .ip(n5522), .ck(clk), .q(
        \cache_data_B[6][70] ) );
  dp_1 \cache_data_B_reg[6][71]  ( .ip(n5521), .ck(clk), .q(
        \cache_data_B[6][71] ) );
  dp_1 \cache_data_B_reg[6][72]  ( .ip(n5520), .ck(clk), .q(
        \cache_data_B[6][72] ) );
  dp_1 \cache_data_B_reg[6][73]  ( .ip(n5519), .ck(clk), .q(
        \cache_data_B[6][73] ) );
  dp_1 \cache_data_B_reg[6][74]  ( .ip(n5518), .ck(clk), .q(
        \cache_data_B[6][74] ) );
  dp_1 \cache_data_B_reg[6][75]  ( .ip(n5517), .ck(clk), .q(
        \cache_data_B[6][75] ) );
  dp_1 \cache_data_B_reg[6][76]  ( .ip(n5516), .ck(clk), .q(
        \cache_data_B[6][76] ) );
  dp_1 \cache_data_B_reg[6][77]  ( .ip(n5515), .ck(clk), .q(
        \cache_data_B[6][77] ) );
  dp_1 \cache_data_B_reg[6][78]  ( .ip(n5514), .ck(clk), .q(
        \cache_data_B[6][78] ) );
  dp_1 \cache_data_B_reg[6][79]  ( .ip(n5513), .ck(clk), .q(
        \cache_data_B[6][79] ) );
  dp_1 \cache_data_B_reg[6][80]  ( .ip(n5512), .ck(clk), .q(
        \cache_data_B[6][80] ) );
  dp_1 \cache_data_B_reg[6][81]  ( .ip(n5511), .ck(clk), .q(
        \cache_data_B[6][81] ) );
  dp_1 \cache_data_B_reg[6][82]  ( .ip(n5510), .ck(clk), .q(
        \cache_data_B[6][82] ) );
  dp_1 \cache_data_B_reg[6][83]  ( .ip(n5509), .ck(clk), .q(
        \cache_data_B[6][83] ) );
  dp_1 \cache_data_B_reg[6][84]  ( .ip(n5508), .ck(clk), .q(
        \cache_data_B[6][84] ) );
  dp_1 \cache_data_B_reg[6][85]  ( .ip(n5507), .ck(clk), .q(
        \cache_data_B[6][85] ) );
  dp_1 \cache_data_B_reg[6][86]  ( .ip(n5506), .ck(clk), .q(
        \cache_data_B[6][86] ) );
  dp_1 \cache_data_B_reg[6][87]  ( .ip(n5505), .ck(clk), .q(
        \cache_data_B[6][87] ) );
  dp_1 \cache_data_B_reg[6][88]  ( .ip(n5504), .ck(clk), .q(
        \cache_data_B[6][88] ) );
  dp_1 \cache_data_B_reg[6][89]  ( .ip(n5503), .ck(clk), .q(
        \cache_data_B[6][89] ) );
  dp_1 \cache_data_B_reg[6][90]  ( .ip(n5502), .ck(clk), .q(
        \cache_data_B[6][90] ) );
  dp_1 \cache_data_B_reg[6][91]  ( .ip(n5501), .ck(clk), .q(
        \cache_data_B[6][91] ) );
  dp_1 \cache_data_B_reg[6][92]  ( .ip(n5500), .ck(clk), .q(
        \cache_data_B[6][92] ) );
  dp_1 \cache_data_B_reg[6][93]  ( .ip(n5499), .ck(clk), .q(
        \cache_data_B[6][93] ) );
  dp_1 \cache_data_B_reg[6][94]  ( .ip(n5498), .ck(clk), .q(
        \cache_data_B[6][94] ) );
  dp_1 \cache_data_B_reg[6][95]  ( .ip(n5497), .ck(clk), .q(
        \cache_data_B[6][95] ) );
  dp_1 \cache_data_B_reg[7][83]  ( .ip(n5400), .ck(clk), .q(
        \cache_data_B[7][83] ) );
  dp_1 \cache_data_B_reg[7][84]  ( .ip(n5399), .ck(clk), .q(
        \cache_data_B[7][84] ) );
  dp_1 \cache_data_B_reg[7][85]  ( .ip(n5398), .ck(clk), .q(
        \cache_data_B[7][85] ) );
  dp_1 \cache_data_B_reg[7][86]  ( .ip(n5397), .ck(clk), .q(
        \cache_data_B[7][86] ) );
  dp_1 \cache_data_B_reg[7][87]  ( .ip(n5396), .ck(clk), .q(
        \cache_data_B[7][87] ) );
  dp_1 \cache_data_B_reg[7][88]  ( .ip(n5395), .ck(clk), .q(
        \cache_data_B[7][88] ) );
  dp_1 \cache_data_B_reg[7][89]  ( .ip(n5394), .ck(clk), .q(
        \cache_data_B[7][89] ) );
  dp_1 \cache_data_B_reg[7][90]  ( .ip(n5393), .ck(clk), .q(
        \cache_data_B[7][90] ) );
  dp_1 \cache_data_B_reg[7][91]  ( .ip(n5392), .ck(clk), .q(
        \cache_data_B[7][91] ) );
  dp_1 \cache_data_B_reg[7][92]  ( .ip(n5391), .ck(clk), .q(
        \cache_data_B[7][92] ) );
  dp_1 \cache_data_B_reg[7][93]  ( .ip(n5390), .ck(clk), .q(
        \cache_data_B[7][93] ) );
  dp_1 \cache_data_B_reg[7][94]  ( .ip(n5389), .ck(clk), .q(
        \cache_data_B[7][94] ) );
  dp_1 \cache_data_B_reg[7][95]  ( .ip(n5388), .ck(clk), .q(
        \cache_data_B[7][95] ) );
  dp_1 \cache_data_B_reg[7][64]  ( .ip(n5387), .ck(clk), .q(
        \cache_data_B[7][64] ) );
  dp_1 \cache_data_B_reg[7][65]  ( .ip(n5386), .ck(clk), .q(
        \cache_data_B[7][65] ) );
  dp_1 \cache_data_B_reg[7][66]  ( .ip(n5385), .ck(clk), .q(
        \cache_data_B[7][66] ) );
  dp_1 \cache_data_B_reg[7][67]  ( .ip(n5384), .ck(clk), .q(
        \cache_data_B[7][67] ) );
  dp_1 \cache_data_B_reg[7][68]  ( .ip(n5383), .ck(clk), .q(
        \cache_data_B[7][68] ) );
  dp_1 \cache_data_B_reg[7][69]  ( .ip(n5382), .ck(clk), .q(
        \cache_data_B[7][69] ) );
  dp_1 \cache_data_B_reg[7][70]  ( .ip(n5381), .ck(clk), .q(
        \cache_data_B[7][70] ) );
  dp_1 \cache_data_B_reg[7][71]  ( .ip(n5380), .ck(clk), .q(
        \cache_data_B[7][71] ) );
  dp_1 \cache_data_B_reg[7][72]  ( .ip(n5379), .ck(clk), .q(
        \cache_data_B[7][72] ) );
  dp_1 \cache_data_B_reg[7][73]  ( .ip(n5378), .ck(clk), .q(
        \cache_data_B[7][73] ) );
  dp_1 \cache_data_B_reg[7][74]  ( .ip(n5377), .ck(clk), .q(
        \cache_data_B[7][74] ) );
  dp_1 \cache_data_B_reg[7][75]  ( .ip(n5376), .ck(clk), .q(
        \cache_data_B[7][75] ) );
  dp_1 \cache_data_B_reg[7][76]  ( .ip(n5375), .ck(clk), .q(
        \cache_data_B[7][76] ) );
  dp_1 \cache_data_B_reg[7][77]  ( .ip(n5374), .ck(clk), .q(
        \cache_data_B[7][77] ) );
  dp_1 \cache_data_B_reg[7][78]  ( .ip(n5373), .ck(clk), .q(
        \cache_data_B[7][78] ) );
  dp_1 \cache_data_B_reg[7][79]  ( .ip(n5372), .ck(clk), .q(
        \cache_data_B[7][79] ) );
  dp_1 \cache_data_B_reg[7][80]  ( .ip(n5371), .ck(clk), .q(
        \cache_data_B[7][80] ) );
  dp_1 \cache_data_B_reg[7][81]  ( .ip(n5370), .ck(clk), .q(
        \cache_data_B[7][81] ) );
  dp_1 \cache_data_B_reg[7][82]  ( .ip(n5369), .ck(clk), .q(
        \cache_data_B[7][82] ) );
  dp_1 \cache_data_B_reg[0][96]  ( .ip(n6264), .ck(clk), .q(
        \cache_data_B[0][96] ) );
  dp_1 \cache_data_B_reg[0][97]  ( .ip(n6263), .ck(clk), .q(
        \cache_data_B[0][97] ) );
  dp_1 \cache_data_B_reg[0][98]  ( .ip(n6262), .ck(clk), .q(
        \cache_data_B[0][98] ) );
  dp_1 \cache_data_B_reg[0][99]  ( .ip(n6261), .ck(clk), .q(
        \cache_data_B[0][99] ) );
  dp_1 \cache_data_B_reg[0][100]  ( .ip(n6260), .ck(clk), .q(
        \cache_data_B[0][100] ) );
  dp_1 \cache_data_B_reg[0][101]  ( .ip(n6259), .ck(clk), .q(
        \cache_data_B[0][101] ) );
  dp_1 \cache_data_B_reg[0][102]  ( .ip(n6258), .ck(clk), .q(
        \cache_data_B[0][102] ) );
  dp_1 \cache_data_B_reg[0][103]  ( .ip(n6257), .ck(clk), .q(
        \cache_data_B[0][103] ) );
  dp_1 \cache_data_B_reg[0][104]  ( .ip(n6256), .ck(clk), .q(
        \cache_data_B[0][104] ) );
  dp_1 \cache_data_B_reg[0][105]  ( .ip(n6255), .ck(clk), .q(
        \cache_data_B[0][105] ) );
  dp_1 \cache_data_B_reg[0][106]  ( .ip(n6254), .ck(clk), .q(
        \cache_data_B[0][106] ) );
  dp_1 \cache_data_B_reg[0][107]  ( .ip(n6253), .ck(clk), .q(
        \cache_data_B[0][107] ) );
  dp_1 \cache_data_B_reg[0][108]  ( .ip(n6252), .ck(clk), .q(
        \cache_data_B[0][108] ) );
  dp_1 \cache_data_B_reg[0][109]  ( .ip(n6251), .ck(clk), .q(
        \cache_data_B[0][109] ) );
  dp_1 \cache_data_B_reg[0][110]  ( .ip(n6250), .ck(clk), .q(
        \cache_data_B[0][110] ) );
  dp_1 \cache_data_B_reg[0][111]  ( .ip(n6249), .ck(clk), .q(
        \cache_data_B[0][111] ) );
  dp_1 \cache_data_B_reg[0][112]  ( .ip(n6248), .ck(clk), .q(
        \cache_data_B[0][112] ) );
  dp_1 \cache_data_B_reg[0][113]  ( .ip(n6247), .ck(clk), .q(
        \cache_data_B[0][113] ) );
  dp_1 \cache_data_B_reg[0][114]  ( .ip(n6246), .ck(clk), .q(
        \cache_data_B[0][114] ) );
  dp_1 \cache_data_B_reg[0][115]  ( .ip(n6245), .ck(clk), .q(
        \cache_data_B[0][115] ) );
  dp_1 \cache_data_B_reg[0][116]  ( .ip(n6244), .ck(clk), .q(
        \cache_data_B[0][116] ) );
  dp_1 \cache_data_B_reg[0][117]  ( .ip(n6243), .ck(clk), .q(
        \cache_data_B[0][117] ) );
  dp_1 \cache_data_B_reg[0][118]  ( .ip(n6242), .ck(clk), .q(
        \cache_data_B[0][118] ) );
  dp_1 \cache_data_B_reg[0][119]  ( .ip(n6241), .ck(clk), .q(
        \cache_data_B[0][119] ) );
  dp_1 \cache_data_B_reg[0][120]  ( .ip(n6240), .ck(clk), .q(
        \cache_data_B[0][120] ) );
  dp_1 \cache_data_B_reg[0][121]  ( .ip(n6239), .ck(clk), .q(
        \cache_data_B[0][121] ) );
  dp_1 \cache_data_B_reg[0][122]  ( .ip(n6238), .ck(clk), .q(
        \cache_data_B[0][122] ) );
  dp_1 \cache_data_B_reg[0][123]  ( .ip(n6237), .ck(clk), .q(
        \cache_data_B[0][123] ) );
  dp_1 \cache_data_B_reg[0][124]  ( .ip(n6236), .ck(clk), .q(
        \cache_data_B[0][124] ) );
  dp_1 \cache_data_B_reg[0][125]  ( .ip(n6235), .ck(clk), .q(
        \cache_data_B[0][125] ) );
  dp_1 \cache_data_B_reg[0][126]  ( .ip(n6234), .ck(clk), .q(
        \cache_data_B[0][126] ) );
  dp_1 \cache_data_B_reg[0][127]  ( .ip(n6233), .ck(clk), .q(
        \cache_data_B[0][127] ) );
  dp_1 \cache_data_B_reg[1][96]  ( .ip(n6136), .ck(clk), .q(
        \cache_data_B[1][96] ) );
  dp_1 \cache_data_B_reg[1][97]  ( .ip(n6135), .ck(clk), .q(
        \cache_data_B[1][97] ) );
  dp_1 \cache_data_B_reg[1][98]  ( .ip(n6134), .ck(clk), .q(
        \cache_data_B[1][98] ) );
  dp_1 \cache_data_B_reg[1][99]  ( .ip(n6133), .ck(clk), .q(
        \cache_data_B[1][99] ) );
  dp_1 \cache_data_B_reg[1][100]  ( .ip(n6132), .ck(clk), .q(
        \cache_data_B[1][100] ) );
  dp_1 \cache_data_B_reg[1][101]  ( .ip(n6131), .ck(clk), .q(
        \cache_data_B[1][101] ) );
  dp_1 \cache_data_B_reg[1][102]  ( .ip(n6130), .ck(clk), .q(
        \cache_data_B[1][102] ) );
  dp_1 \cache_data_B_reg[1][103]  ( .ip(n6129), .ck(clk), .q(
        \cache_data_B[1][103] ) );
  dp_1 \cache_data_B_reg[1][104]  ( .ip(n6128), .ck(clk), .q(
        \cache_data_B[1][104] ) );
  dp_1 \cache_data_B_reg[1][105]  ( .ip(n6127), .ck(clk), .q(
        \cache_data_B[1][105] ) );
  dp_1 \cache_data_B_reg[1][106]  ( .ip(n6126), .ck(clk), .q(
        \cache_data_B[1][106] ) );
  dp_1 \cache_data_B_reg[1][107]  ( .ip(n6125), .ck(clk), .q(
        \cache_data_B[1][107] ) );
  dp_1 \cache_data_B_reg[1][108]  ( .ip(n6124), .ck(clk), .q(
        \cache_data_B[1][108] ) );
  dp_1 \cache_data_B_reg[1][109]  ( .ip(n6123), .ck(clk), .q(
        \cache_data_B[1][109] ) );
  dp_1 \cache_data_B_reg[1][110]  ( .ip(n6122), .ck(clk), .q(
        \cache_data_B[1][110] ) );
  dp_1 \cache_data_B_reg[1][111]  ( .ip(n6121), .ck(clk), .q(
        \cache_data_B[1][111] ) );
  dp_1 \cache_data_B_reg[1][112]  ( .ip(n6120), .ck(clk), .q(
        \cache_data_B[1][112] ) );
  dp_1 \cache_data_B_reg[1][113]  ( .ip(n6119), .ck(clk), .q(
        \cache_data_B[1][113] ) );
  dp_1 \cache_data_B_reg[1][114]  ( .ip(n6118), .ck(clk), .q(
        \cache_data_B[1][114] ) );
  dp_1 \cache_data_B_reg[1][115]  ( .ip(n6117), .ck(clk), .q(
        \cache_data_B[1][115] ) );
  dp_1 \cache_data_B_reg[1][116]  ( .ip(n6116), .ck(clk), .q(
        \cache_data_B[1][116] ) );
  dp_1 \cache_data_B_reg[1][117]  ( .ip(n6115), .ck(clk), .q(
        \cache_data_B[1][117] ) );
  dp_1 \cache_data_B_reg[1][118]  ( .ip(n6114), .ck(clk), .q(
        \cache_data_B[1][118] ) );
  dp_1 \cache_data_B_reg[1][119]  ( .ip(n6113), .ck(clk), .q(
        \cache_data_B[1][119] ) );
  dp_1 \cache_data_B_reg[1][120]  ( .ip(n6112), .ck(clk), .q(
        \cache_data_B[1][120] ) );
  dp_1 \cache_data_B_reg[1][121]  ( .ip(n6111), .ck(clk), .q(
        \cache_data_B[1][121] ) );
  dp_1 \cache_data_B_reg[1][122]  ( .ip(n6110), .ck(clk), .q(
        \cache_data_B[1][122] ) );
  dp_1 \cache_data_B_reg[1][123]  ( .ip(n6109), .ck(clk), .q(
        \cache_data_B[1][123] ) );
  dp_1 \cache_data_B_reg[1][124]  ( .ip(n6108), .ck(clk), .q(
        \cache_data_B[1][124] ) );
  dp_1 \cache_data_B_reg[1][125]  ( .ip(n6107), .ck(clk), .q(
        \cache_data_B[1][125] ) );
  dp_1 \cache_data_B_reg[1][126]  ( .ip(n6106), .ck(clk), .q(
        \cache_data_B[1][126] ) );
  dp_1 \cache_data_B_reg[1][127]  ( .ip(n6105), .ck(clk), .q(
        \cache_data_B[1][127] ) );
  dp_1 \cache_data_B_reg[2][96]  ( .ip(n6008), .ck(clk), .q(
        \cache_data_B[2][96] ) );
  dp_1 \cache_data_B_reg[2][97]  ( .ip(n6007), .ck(clk), .q(
        \cache_data_B[2][97] ) );
  dp_1 \cache_data_B_reg[2][98]  ( .ip(n6006), .ck(clk), .q(
        \cache_data_B[2][98] ) );
  dp_1 \cache_data_B_reg[2][99]  ( .ip(n6005), .ck(clk), .q(
        \cache_data_B[2][99] ) );
  dp_1 \cache_data_B_reg[2][100]  ( .ip(n6004), .ck(clk), .q(
        \cache_data_B[2][100] ) );
  dp_1 \cache_data_B_reg[2][101]  ( .ip(n6003), .ck(clk), .q(
        \cache_data_B[2][101] ) );
  dp_1 \cache_data_B_reg[2][102]  ( .ip(n6002), .ck(clk), .q(
        \cache_data_B[2][102] ) );
  dp_1 \cache_data_B_reg[2][103]  ( .ip(n6001), .ck(clk), .q(
        \cache_data_B[2][103] ) );
  dp_1 \cache_data_B_reg[2][104]  ( .ip(n6000), .ck(clk), .q(
        \cache_data_B[2][104] ) );
  dp_1 \cache_data_B_reg[2][105]  ( .ip(n5999), .ck(clk), .q(
        \cache_data_B[2][105] ) );
  dp_1 \cache_data_B_reg[2][106]  ( .ip(n5998), .ck(clk), .q(
        \cache_data_B[2][106] ) );
  dp_1 \cache_data_B_reg[2][107]  ( .ip(n5997), .ck(clk), .q(
        \cache_data_B[2][107] ) );
  dp_1 \cache_data_B_reg[2][108]  ( .ip(n5996), .ck(clk), .q(
        \cache_data_B[2][108] ) );
  dp_1 \cache_data_B_reg[2][109]  ( .ip(n5995), .ck(clk), .q(
        \cache_data_B[2][109] ) );
  dp_1 \cache_data_B_reg[2][110]  ( .ip(n5994), .ck(clk), .q(
        \cache_data_B[2][110] ) );
  dp_1 \cache_data_B_reg[2][111]  ( .ip(n5993), .ck(clk), .q(
        \cache_data_B[2][111] ) );
  dp_1 \cache_data_B_reg[2][112]  ( .ip(n5992), .ck(clk), .q(
        \cache_data_B[2][112] ) );
  dp_1 \cache_data_B_reg[2][113]  ( .ip(n5991), .ck(clk), .q(
        \cache_data_B[2][113] ) );
  dp_1 \cache_data_B_reg[2][114]  ( .ip(n5990), .ck(clk), .q(
        \cache_data_B[2][114] ) );
  dp_1 \cache_data_B_reg[2][115]  ( .ip(n5989), .ck(clk), .q(
        \cache_data_B[2][115] ) );
  dp_1 \cache_data_B_reg[2][116]  ( .ip(n5988), .ck(clk), .q(
        \cache_data_B[2][116] ) );
  dp_1 \cache_data_B_reg[2][117]  ( .ip(n5987), .ck(clk), .q(
        \cache_data_B[2][117] ) );
  dp_1 \cache_data_B_reg[2][118]  ( .ip(n5986), .ck(clk), .q(
        \cache_data_B[2][118] ) );
  dp_1 \cache_data_B_reg[2][119]  ( .ip(n5985), .ck(clk), .q(
        \cache_data_B[2][119] ) );
  dp_1 \cache_data_B_reg[2][120]  ( .ip(n5984), .ck(clk), .q(
        \cache_data_B[2][120] ) );
  dp_1 \cache_data_B_reg[2][121]  ( .ip(n5983), .ck(clk), .q(
        \cache_data_B[2][121] ) );
  dp_1 \cache_data_B_reg[2][122]  ( .ip(n5982), .ck(clk), .q(
        \cache_data_B[2][122] ) );
  dp_1 \cache_data_B_reg[2][123]  ( .ip(n5981), .ck(clk), .q(
        \cache_data_B[2][123] ) );
  dp_1 \cache_data_B_reg[2][124]  ( .ip(n5980), .ck(clk), .q(
        \cache_data_B[2][124] ) );
  dp_1 \cache_data_B_reg[2][125]  ( .ip(n5979), .ck(clk), .q(
        \cache_data_B[2][125] ) );
  dp_1 \cache_data_B_reg[2][126]  ( .ip(n5978), .ck(clk), .q(
        \cache_data_B[2][126] ) );
  dp_1 \cache_data_B_reg[2][127]  ( .ip(n5977), .ck(clk), .q(
        \cache_data_B[2][127] ) );
  dp_1 \cache_data_B_reg[3][100]  ( .ip(n5880), .ck(clk), .q(
        \cache_data_B[3][100] ) );
  dp_1 \cache_data_B_reg[3][101]  ( .ip(n5879), .ck(clk), .q(
        \cache_data_B[3][101] ) );
  dp_1 \cache_data_B_reg[3][102]  ( .ip(n5878), .ck(clk), .q(
        \cache_data_B[3][102] ) );
  dp_1 \cache_data_B_reg[3][103]  ( .ip(n5877), .ck(clk), .q(
        \cache_data_B[3][103] ) );
  dp_1 \cache_data_B_reg[3][104]  ( .ip(n5876), .ck(clk), .q(
        \cache_data_B[3][104] ) );
  dp_1 \cache_data_B_reg[3][105]  ( .ip(n5875), .ck(clk), .q(
        \cache_data_B[3][105] ) );
  dp_1 \cache_data_B_reg[3][106]  ( .ip(n5874), .ck(clk), .q(
        \cache_data_B[3][106] ) );
  dp_1 \cache_data_B_reg[3][107]  ( .ip(n5873), .ck(clk), .q(
        \cache_data_B[3][107] ) );
  dp_1 \cache_data_B_reg[3][108]  ( .ip(n5872), .ck(clk), .q(
        \cache_data_B[3][108] ) );
  dp_1 \cache_data_B_reg[3][109]  ( .ip(n5871), .ck(clk), .q(
        \cache_data_B[3][109] ) );
  dp_1 \cache_data_B_reg[3][110]  ( .ip(n5870), .ck(clk), .q(
        \cache_data_B[3][110] ) );
  dp_1 \cache_data_B_reg[3][111]  ( .ip(n5869), .ck(clk), .q(
        \cache_data_B[3][111] ) );
  dp_1 \cache_data_B_reg[3][112]  ( .ip(n5868), .ck(clk), .q(
        \cache_data_B[3][112] ) );
  dp_1 \cache_data_B_reg[3][113]  ( .ip(n5867), .ck(clk), .q(
        \cache_data_B[3][113] ) );
  dp_1 \cache_data_B_reg[3][114]  ( .ip(n5866), .ck(clk), .q(
        \cache_data_B[3][114] ) );
  dp_1 \cache_data_B_reg[3][115]  ( .ip(n5865), .ck(clk), .q(
        \cache_data_B[3][115] ) );
  dp_1 \cache_data_B_reg[3][116]  ( .ip(n5864), .ck(clk), .q(
        \cache_data_B[3][116] ) );
  dp_1 \cache_data_B_reg[3][117]  ( .ip(n5863), .ck(clk), .q(
        \cache_data_B[3][117] ) );
  dp_1 \cache_data_B_reg[3][118]  ( .ip(n5862), .ck(clk), .q(
        \cache_data_B[3][118] ) );
  dp_1 \cache_data_B_reg[3][119]  ( .ip(n5861), .ck(clk), .q(
        \cache_data_B[3][119] ) );
  dp_1 \cache_data_B_reg[3][120]  ( .ip(n5860), .ck(clk), .q(
        \cache_data_B[3][120] ) );
  dp_1 \cache_data_B_reg[3][121]  ( .ip(n5859), .ck(clk), .q(
        \cache_data_B[3][121] ) );
  dp_1 \cache_data_B_reg[3][122]  ( .ip(n5858), .ck(clk), .q(
        \cache_data_B[3][122] ) );
  dp_1 \cache_data_B_reg[3][123]  ( .ip(n5857), .ck(clk), .q(
        \cache_data_B[3][123] ) );
  dp_1 \cache_data_B_reg[3][124]  ( .ip(n5856), .ck(clk), .q(
        \cache_data_B[3][124] ) );
  dp_1 \cache_data_B_reg[3][125]  ( .ip(n5855), .ck(clk), .q(
        \cache_data_B[3][125] ) );
  dp_1 \cache_data_B_reg[3][126]  ( .ip(n5854), .ck(clk), .q(
        \cache_data_B[3][126] ) );
  dp_1 \cache_data_B_reg[3][127]  ( .ip(n5853), .ck(clk), .q(
        \cache_data_B[3][127] ) );
  dp_1 \cache_data_B_reg[3][96]  ( .ip(n5852), .ck(clk), .q(
        \cache_data_B[3][96] ) );
  dp_1 \cache_data_B_reg[3][97]  ( .ip(n5851), .ck(clk), .q(
        \cache_data_B[3][97] ) );
  dp_1 \cache_data_B_reg[3][98]  ( .ip(n5850), .ck(clk), .q(
        \cache_data_B[3][98] ) );
  dp_1 \cache_data_B_reg[3][99]  ( .ip(n5849), .ck(clk), .q(
        \cache_data_B[3][99] ) );
  dp_1 \cache_data_B_reg[4][96]  ( .ip(n5752), .ck(clk), .q(
        \cache_data_B[4][96] ) );
  dp_1 \cache_data_B_reg[4][97]  ( .ip(n5751), .ck(clk), .q(
        \cache_data_B[4][97] ) );
  dp_1 \cache_data_B_reg[4][98]  ( .ip(n5750), .ck(clk), .q(
        \cache_data_B[4][98] ) );
  dp_1 \cache_data_B_reg[4][99]  ( .ip(n5749), .ck(clk), .q(
        \cache_data_B[4][99] ) );
  dp_1 \cache_data_B_reg[4][100]  ( .ip(n5748), .ck(clk), .q(
        \cache_data_B[4][100] ) );
  dp_1 \cache_data_B_reg[4][101]  ( .ip(n5747), .ck(clk), .q(
        \cache_data_B[4][101] ) );
  dp_1 \cache_data_B_reg[4][102]  ( .ip(n5746), .ck(clk), .q(
        \cache_data_B[4][102] ) );
  dp_1 \cache_data_B_reg[4][103]  ( .ip(n5745), .ck(clk), .q(
        \cache_data_B[4][103] ) );
  dp_1 \cache_data_B_reg[4][104]  ( .ip(n5744), .ck(clk), .q(
        \cache_data_B[4][104] ) );
  dp_1 \cache_data_B_reg[4][105]  ( .ip(n5743), .ck(clk), .q(
        \cache_data_B[4][105] ) );
  dp_1 \cache_data_B_reg[4][106]  ( .ip(n5742), .ck(clk), .q(
        \cache_data_B[4][106] ) );
  dp_1 \cache_data_B_reg[4][107]  ( .ip(n5741), .ck(clk), .q(
        \cache_data_B[4][107] ) );
  dp_1 \cache_data_B_reg[4][108]  ( .ip(n5740), .ck(clk), .q(
        \cache_data_B[4][108] ) );
  dp_1 \cache_data_B_reg[4][109]  ( .ip(n5739), .ck(clk), .q(
        \cache_data_B[4][109] ) );
  dp_1 \cache_data_B_reg[4][110]  ( .ip(n5738), .ck(clk), .q(
        \cache_data_B[4][110] ) );
  dp_1 \cache_data_B_reg[4][111]  ( .ip(n5737), .ck(clk), .q(
        \cache_data_B[4][111] ) );
  dp_1 \cache_data_B_reg[4][112]  ( .ip(n5736), .ck(clk), .q(
        \cache_data_B[4][112] ) );
  dp_1 \cache_data_B_reg[4][113]  ( .ip(n5735), .ck(clk), .q(
        \cache_data_B[4][113] ) );
  dp_1 \cache_data_B_reg[4][114]  ( .ip(n5734), .ck(clk), .q(
        \cache_data_B[4][114] ) );
  dp_1 \cache_data_B_reg[4][115]  ( .ip(n5733), .ck(clk), .q(
        \cache_data_B[4][115] ) );
  dp_1 \cache_data_B_reg[4][116]  ( .ip(n5732), .ck(clk), .q(
        \cache_data_B[4][116] ) );
  dp_1 \cache_data_B_reg[4][117]  ( .ip(n5731), .ck(clk), .q(
        \cache_data_B[4][117] ) );
  dp_1 \cache_data_B_reg[4][118]  ( .ip(n5730), .ck(clk), .q(
        \cache_data_B[4][118] ) );
  dp_1 \cache_data_B_reg[4][119]  ( .ip(n5729), .ck(clk), .q(
        \cache_data_B[4][119] ) );
  dp_1 \cache_data_B_reg[4][120]  ( .ip(n5728), .ck(clk), .q(
        \cache_data_B[4][120] ) );
  dp_1 \cache_data_B_reg[4][121]  ( .ip(n5727), .ck(clk), .q(
        \cache_data_B[4][121] ) );
  dp_1 \cache_data_B_reg[4][122]  ( .ip(n5726), .ck(clk), .q(
        \cache_data_B[4][122] ) );
  dp_1 \cache_data_B_reg[4][123]  ( .ip(n5725), .ck(clk), .q(
        \cache_data_B[4][123] ) );
  dp_1 \cache_data_B_reg[4][124]  ( .ip(n5724), .ck(clk), .q(
        \cache_data_B[4][124] ) );
  dp_1 \cache_data_B_reg[4][125]  ( .ip(n5723), .ck(clk), .q(
        \cache_data_B[4][125] ) );
  dp_1 \cache_data_B_reg[4][126]  ( .ip(n5722), .ck(clk), .q(
        \cache_data_B[4][126] ) );
  dp_1 \cache_data_B_reg[4][127]  ( .ip(n5721), .ck(clk), .q(
        \cache_data_B[4][127] ) );
  dp_1 \cache_data_B_reg[5][96]  ( .ip(n5624), .ck(clk), .q(
        \cache_data_B[5][96] ) );
  dp_1 \cache_data_B_reg[5][97]  ( .ip(n5623), .ck(clk), .q(
        \cache_data_B[5][97] ) );
  dp_1 \cache_data_B_reg[5][98]  ( .ip(n5622), .ck(clk), .q(
        \cache_data_B[5][98] ) );
  dp_1 \cache_data_B_reg[5][99]  ( .ip(n5621), .ck(clk), .q(
        \cache_data_B[5][99] ) );
  dp_1 \cache_data_B_reg[5][100]  ( .ip(n5620), .ck(clk), .q(
        \cache_data_B[5][100] ) );
  dp_1 \cache_data_B_reg[5][101]  ( .ip(n5619), .ck(clk), .q(
        \cache_data_B[5][101] ) );
  dp_1 \cache_data_B_reg[5][102]  ( .ip(n5618), .ck(clk), .q(
        \cache_data_B[5][102] ) );
  dp_1 \cache_data_B_reg[5][103]  ( .ip(n5617), .ck(clk), .q(
        \cache_data_B[5][103] ) );
  dp_1 \cache_data_B_reg[5][104]  ( .ip(n5616), .ck(clk), .q(
        \cache_data_B[5][104] ) );
  dp_1 \cache_data_B_reg[5][105]  ( .ip(n5615), .ck(clk), .q(
        \cache_data_B[5][105] ) );
  dp_1 \cache_data_B_reg[5][106]  ( .ip(n5614), .ck(clk), .q(
        \cache_data_B[5][106] ) );
  dp_1 \cache_data_B_reg[5][107]  ( .ip(n5613), .ck(clk), .q(
        \cache_data_B[5][107] ) );
  dp_1 \cache_data_B_reg[5][108]  ( .ip(n5612), .ck(clk), .q(
        \cache_data_B[5][108] ) );
  dp_1 \cache_data_B_reg[5][109]  ( .ip(n5611), .ck(clk), .q(
        \cache_data_B[5][109] ) );
  dp_1 \cache_data_B_reg[5][110]  ( .ip(n5610), .ck(clk), .q(
        \cache_data_B[5][110] ) );
  dp_1 \cache_data_B_reg[5][111]  ( .ip(n5609), .ck(clk), .q(
        \cache_data_B[5][111] ) );
  dp_1 \cache_data_B_reg[5][112]  ( .ip(n5608), .ck(clk), .q(
        \cache_data_B[5][112] ) );
  dp_1 \cache_data_B_reg[5][113]  ( .ip(n5607), .ck(clk), .q(
        \cache_data_B[5][113] ) );
  dp_1 \cache_data_B_reg[5][114]  ( .ip(n5606), .ck(clk), .q(
        \cache_data_B[5][114] ) );
  dp_1 \cache_data_B_reg[5][115]  ( .ip(n5605), .ck(clk), .q(
        \cache_data_B[5][115] ) );
  dp_1 \cache_data_B_reg[5][116]  ( .ip(n5604), .ck(clk), .q(
        \cache_data_B[5][116] ) );
  dp_1 \cache_data_B_reg[5][117]  ( .ip(n5603), .ck(clk), .q(
        \cache_data_B[5][117] ) );
  dp_1 \cache_data_B_reg[5][118]  ( .ip(n5602), .ck(clk), .q(
        \cache_data_B[5][118] ) );
  dp_1 \cache_data_B_reg[5][119]  ( .ip(n5601), .ck(clk), .q(
        \cache_data_B[5][119] ) );
  dp_1 \cache_data_B_reg[5][120]  ( .ip(n5600), .ck(clk), .q(
        \cache_data_B[5][120] ) );
  dp_1 \cache_data_B_reg[5][121]  ( .ip(n5599), .ck(clk), .q(
        \cache_data_B[5][121] ) );
  dp_1 \cache_data_B_reg[5][122]  ( .ip(n5598), .ck(clk), .q(
        \cache_data_B[5][122] ) );
  dp_1 \cache_data_B_reg[5][123]  ( .ip(n5597), .ck(clk), .q(
        \cache_data_B[5][123] ) );
  dp_1 \cache_data_B_reg[5][124]  ( .ip(n5596), .ck(clk), .q(
        \cache_data_B[5][124] ) );
  dp_1 \cache_data_B_reg[5][125]  ( .ip(n5595), .ck(clk), .q(
        \cache_data_B[5][125] ) );
  dp_1 \cache_data_B_reg[5][126]  ( .ip(n5594), .ck(clk), .q(
        \cache_data_B[5][126] ) );
  dp_1 \cache_data_B_reg[5][127]  ( .ip(n5593), .ck(clk), .q(
        \cache_data_B[5][127] ) );
  dp_1 \cache_data_B_reg[6][112]  ( .ip(n5496), .ck(clk), .q(
        \cache_data_B[6][112] ) );
  dp_1 \cache_data_B_reg[6][113]  ( .ip(n5495), .ck(clk), .q(
        \cache_data_B[6][113] ) );
  dp_1 \cache_data_B_reg[6][114]  ( .ip(n5494), .ck(clk), .q(
        \cache_data_B[6][114] ) );
  dp_1 \cache_data_B_reg[6][115]  ( .ip(n5493), .ck(clk), .q(
        \cache_data_B[6][115] ) );
  dp_1 \cache_data_B_reg[6][116]  ( .ip(n5492), .ck(clk), .q(
        \cache_data_B[6][116] ) );
  dp_1 \cache_data_B_reg[6][117]  ( .ip(n5491), .ck(clk), .q(
        \cache_data_B[6][117] ) );
  dp_1 \cache_data_B_reg[6][118]  ( .ip(n5490), .ck(clk), .q(
        \cache_data_B[6][118] ) );
  dp_1 \cache_data_B_reg[6][119]  ( .ip(n5489), .ck(clk), .q(
        \cache_data_B[6][119] ) );
  dp_1 \cache_data_B_reg[6][120]  ( .ip(n5488), .ck(clk), .q(
        \cache_data_B[6][120] ) );
  dp_1 \cache_data_B_reg[6][121]  ( .ip(n5487), .ck(clk), .q(
        \cache_data_B[6][121] ) );
  dp_1 \cache_data_B_reg[6][122]  ( .ip(n5486), .ck(clk), .q(
        \cache_data_B[6][122] ) );
  dp_1 \cache_data_B_reg[6][123]  ( .ip(n5485), .ck(clk), .q(
        \cache_data_B[6][123] ) );
  dp_1 \cache_data_B_reg[6][124]  ( .ip(n5484), .ck(clk), .q(
        \cache_data_B[6][124] ) );
  dp_1 \cache_data_B_reg[6][125]  ( .ip(n5483), .ck(clk), .q(
        \cache_data_B[6][125] ) );
  dp_1 \cache_data_B_reg[6][126]  ( .ip(n5482), .ck(clk), .q(
        \cache_data_B[6][126] ) );
  dp_1 \cache_data_B_reg[6][127]  ( .ip(n5481), .ck(clk), .q(
        \cache_data_B[6][127] ) );
  dp_1 \cache_data_B_reg[6][96]  ( .ip(n5480), .ck(clk), .q(
        \cache_data_B[6][96] ) );
  dp_1 \cache_data_B_reg[6][97]  ( .ip(n5479), .ck(clk), .q(
        \cache_data_B[6][97] ) );
  dp_1 \cache_data_B_reg[6][98]  ( .ip(n5478), .ck(clk), .q(
        \cache_data_B[6][98] ) );
  dp_1 \cache_data_B_reg[6][99]  ( .ip(n5477), .ck(clk), .q(
        \cache_data_B[6][99] ) );
  dp_1 \cache_data_B_reg[6][100]  ( .ip(n5476), .ck(clk), .q(
        \cache_data_B[6][100] ) );
  dp_1 \cache_data_B_reg[6][101]  ( .ip(n5475), .ck(clk), .q(
        \cache_data_B[6][101] ) );
  dp_1 \cache_data_B_reg[6][102]  ( .ip(n5474), .ck(clk), .q(
        \cache_data_B[6][102] ) );
  dp_1 \cache_data_B_reg[6][103]  ( .ip(n5473), .ck(clk), .q(
        \cache_data_B[6][103] ) );
  dp_1 \cache_data_B_reg[6][104]  ( .ip(n5472), .ck(clk), .q(
        \cache_data_B[6][104] ) );
  dp_1 \cache_data_B_reg[6][105]  ( .ip(n5471), .ck(clk), .q(
        \cache_data_B[6][105] ) );
  dp_1 \cache_data_B_reg[6][106]  ( .ip(n5470), .ck(clk), .q(
        \cache_data_B[6][106] ) );
  dp_1 \cache_data_B_reg[6][107]  ( .ip(n5469), .ck(clk), .q(
        \cache_data_B[6][107] ) );
  dp_1 \cache_data_B_reg[6][108]  ( .ip(n5468), .ck(clk), .q(
        \cache_data_B[6][108] ) );
  dp_1 \cache_data_B_reg[6][109]  ( .ip(n5467), .ck(clk), .q(
        \cache_data_B[6][109] ) );
  dp_1 \cache_data_B_reg[6][110]  ( .ip(n5466), .ck(clk), .q(
        \cache_data_B[6][110] ) );
  dp_1 \cache_data_B_reg[6][111]  ( .ip(n5465), .ck(clk), .q(
        \cache_data_B[6][111] ) );
  dp_1 \cache_data_B_reg[7][96]  ( .ip(n5368), .ck(clk), .q(
        \cache_data_B[7][96] ) );
  dp_1 \cache_data_B_reg[7][97]  ( .ip(n5367), .ck(clk), .q(
        \cache_data_B[7][97] ) );
  dp_1 \cache_data_B_reg[7][98]  ( .ip(n5366), .ck(clk), .q(
        \cache_data_B[7][98] ) );
  dp_1 \cache_data_B_reg[7][99]  ( .ip(n5365), .ck(clk), .q(
        \cache_data_B[7][99] ) );
  dp_1 \cache_data_B_reg[7][100]  ( .ip(n5364), .ck(clk), .q(
        \cache_data_B[7][100] ) );
  dp_1 \cache_data_B_reg[7][101]  ( .ip(n5363), .ck(clk), .q(
        \cache_data_B[7][101] ) );
  dp_1 \cache_data_B_reg[7][102]  ( .ip(n5362), .ck(clk), .q(
        \cache_data_B[7][102] ) );
  dp_1 \cache_data_B_reg[7][103]  ( .ip(n5361), .ck(clk), .q(
        \cache_data_B[7][103] ) );
  dp_1 \cache_data_B_reg[7][104]  ( .ip(n5360), .ck(clk), .q(
        \cache_data_B[7][104] ) );
  dp_1 \cache_data_B_reg[7][105]  ( .ip(n5359), .ck(clk), .q(
        \cache_data_B[7][105] ) );
  dp_1 \cache_data_B_reg[7][106]  ( .ip(n5358), .ck(clk), .q(
        \cache_data_B[7][106] ) );
  dp_1 \cache_data_B_reg[7][107]  ( .ip(n5357), .ck(clk), .q(
        \cache_data_B[7][107] ) );
  dp_1 \cache_data_B_reg[7][108]  ( .ip(n5356), .ck(clk), .q(
        \cache_data_B[7][108] ) );
  dp_1 \cache_data_B_reg[7][109]  ( .ip(n5355), .ck(clk), .q(
        \cache_data_B[7][109] ) );
  dp_1 \cache_data_B_reg[7][110]  ( .ip(n5354), .ck(clk), .q(
        \cache_data_B[7][110] ) );
  dp_1 \cache_data_B_reg[7][111]  ( .ip(n5353), .ck(clk), .q(
        \cache_data_B[7][111] ) );
  dp_1 \cache_data_B_reg[7][112]  ( .ip(n5352), .ck(clk), .q(
        \cache_data_B[7][112] ) );
  dp_1 \cache_data_B_reg[7][113]  ( .ip(n5351), .ck(clk), .q(
        \cache_data_B[7][113] ) );
  dp_1 \cache_data_B_reg[7][114]  ( .ip(n5350), .ck(clk), .q(
        \cache_data_B[7][114] ) );
  dp_1 \cache_data_B_reg[7][115]  ( .ip(n5349), .ck(clk), .q(
        \cache_data_B[7][115] ) );
  dp_1 \cache_data_B_reg[7][116]  ( .ip(n5348), .ck(clk), .q(
        \cache_data_B[7][116] ) );
  dp_1 \cache_data_B_reg[7][117]  ( .ip(n5347), .ck(clk), .q(
        \cache_data_B[7][117] ) );
  dp_1 \cache_data_B_reg[7][118]  ( .ip(n5346), .ck(clk), .q(
        \cache_data_B[7][118] ) );
  dp_1 \cache_data_B_reg[7][119]  ( .ip(n5345), .ck(clk), .q(
        \cache_data_B[7][119] ) );
  dp_1 \cache_data_B_reg[7][120]  ( .ip(n5344), .ck(clk), .q(
        \cache_data_B[7][120] ) );
  dp_1 \cache_data_B_reg[7][121]  ( .ip(n5343), .ck(clk), .q(
        \cache_data_B[7][121] ) );
  dp_1 \cache_data_B_reg[7][122]  ( .ip(n5342), .ck(clk), .q(
        \cache_data_B[7][122] ) );
  dp_1 \cache_data_B_reg[7][123]  ( .ip(n5341), .ck(clk), .q(
        \cache_data_B[7][123] ) );
  dp_1 \cache_data_B_reg[7][124]  ( .ip(n5340), .ck(clk), .q(
        \cache_data_B[7][124] ) );
  dp_1 \cache_data_B_reg[7][125]  ( .ip(n5339), .ck(clk), .q(
        \cache_data_B[7][125] ) );
  dp_1 \cache_data_B_reg[7][126]  ( .ip(n5338), .ck(clk), .q(
        \cache_data_B[7][126] ) );
  dp_1 \cache_data_B_reg[7][127]  ( .ip(n5337), .ck(clk), .q(
        \cache_data_B[7][127] ) );
  dp_1 \cache_data_A_reg[0][25]  ( .ip(n7384), .ck(clk), .q(
        \cache_data_A[0][25] ) );
  dp_1 \cache_data_A_reg[0][26]  ( .ip(n7383), .ck(clk), .q(
        \cache_data_A[0][26] ) );
  dp_1 \cache_data_A_reg[0][27]  ( .ip(n7382), .ck(clk), .q(
        \cache_data_A[0][27] ) );
  dp_1 \cache_data_A_reg[0][28]  ( .ip(n7381), .ck(clk), .q(
        \cache_data_A[0][28] ) );
  dp_1 \cache_data_A_reg[0][29]  ( .ip(n7380), .ck(clk), .q(
        \cache_data_A[0][29] ) );
  dp_1 \cache_data_A_reg[0][30]  ( .ip(n7379), .ck(clk), .q(
        \cache_data_A[0][30] ) );
  dp_1 \cache_data_A_reg[0][31]  ( .ip(n7378), .ck(clk), .q(
        \cache_data_A[0][31] ) );
  dp_1 \cache_data_A_reg[0][0]  ( .ip(n7377), .ck(clk), .q(
        \cache_data_A[0][0] ) );
  dp_1 \cache_data_A_reg[0][1]  ( .ip(n7376), .ck(clk), .q(
        \cache_data_A[0][1] ) );
  dp_1 \cache_data_A_reg[0][2]  ( .ip(n7375), .ck(clk), .q(
        \cache_data_A[0][2] ) );
  dp_1 \cache_data_A_reg[0][3]  ( .ip(n7374), .ck(clk), .q(
        \cache_data_A[0][3] ) );
  dp_1 \cache_data_A_reg[0][4]  ( .ip(n7373), .ck(clk), .q(
        \cache_data_A[0][4] ) );
  dp_1 \cache_data_A_reg[0][5]  ( .ip(n7372), .ck(clk), .q(
        \cache_data_A[0][5] ) );
  dp_1 \cache_data_A_reg[0][6]  ( .ip(n7371), .ck(clk), .q(
        \cache_data_A[0][6] ) );
  dp_1 \cache_data_A_reg[0][7]  ( .ip(n7370), .ck(clk), .q(
        \cache_data_A[0][7] ) );
  dp_1 \cache_data_A_reg[0][8]  ( .ip(n7369), .ck(clk), .q(
        \cache_data_A[0][8] ) );
  dp_1 \cache_data_A_reg[0][9]  ( .ip(n7368), .ck(clk), .q(
        \cache_data_A[0][9] ) );
  dp_1 \cache_data_A_reg[0][10]  ( .ip(n7367), .ck(clk), .q(
        \cache_data_A[0][10] ) );
  dp_1 \cache_data_A_reg[0][11]  ( .ip(n7366), .ck(clk), .q(
        \cache_data_A[0][11] ) );
  dp_1 \cache_data_A_reg[0][12]  ( .ip(n7365), .ck(clk), .q(
        \cache_data_A[0][12] ) );
  dp_1 \cache_data_A_reg[0][13]  ( .ip(n7364), .ck(clk), .q(
        \cache_data_A[0][13] ) );
  dp_1 \cache_data_A_reg[0][14]  ( .ip(n7363), .ck(clk), .q(
        \cache_data_A[0][14] ) );
  dp_1 \cache_data_A_reg[0][15]  ( .ip(n7362), .ck(clk), .q(
        \cache_data_A[0][15] ) );
  dp_1 \cache_data_A_reg[0][16]  ( .ip(n7361), .ck(clk), .q(
        \cache_data_A[0][16] ) );
  dp_1 \cache_data_A_reg[0][17]  ( .ip(n7360), .ck(clk), .q(
        \cache_data_A[0][17] ) );
  dp_1 \cache_data_A_reg[0][18]  ( .ip(n7359), .ck(clk), .q(
        \cache_data_A[0][18] ) );
  dp_1 \cache_data_A_reg[0][19]  ( .ip(n7358), .ck(clk), .q(
        \cache_data_A[0][19] ) );
  dp_1 \cache_data_A_reg[0][20]  ( .ip(n7357), .ck(clk), .q(
        \cache_data_A[0][20] ) );
  dp_1 \cache_data_A_reg[0][21]  ( .ip(n7356), .ck(clk), .q(
        \cache_data_A[0][21] ) );
  dp_1 \cache_data_A_reg[0][22]  ( .ip(n7355), .ck(clk), .q(
        \cache_data_A[0][22] ) );
  dp_1 \cache_data_A_reg[0][23]  ( .ip(n7354), .ck(clk), .q(
        \cache_data_A[0][23] ) );
  dp_1 \cache_data_A_reg[0][24]  ( .ip(n7353), .ck(clk), .q(
        \cache_data_A[0][24] ) );
  dp_1 \cache_data_A_reg[1][0]  ( .ip(n7256), .ck(clk), .q(
        \cache_data_A[1][0] ) );
  dp_1 \cache_data_A_reg[1][1]  ( .ip(n7255), .ck(clk), .q(
        \cache_data_A[1][1] ) );
  dp_1 \cache_data_A_reg[1][2]  ( .ip(n7254), .ck(clk), .q(
        \cache_data_A[1][2] ) );
  dp_1 \cache_data_A_reg[1][3]  ( .ip(n7253), .ck(clk), .q(
        \cache_data_A[1][3] ) );
  dp_1 \cache_data_A_reg[1][4]  ( .ip(n7252), .ck(clk), .q(
        \cache_data_A[1][4] ) );
  dp_1 \cache_data_A_reg[1][5]  ( .ip(n7251), .ck(clk), .q(
        \cache_data_A[1][5] ) );
  dp_1 \cache_data_A_reg[1][6]  ( .ip(n7250), .ck(clk), .q(
        \cache_data_A[1][6] ) );
  dp_1 \cache_data_A_reg[1][7]  ( .ip(n7249), .ck(clk), .q(
        \cache_data_A[1][7] ) );
  dp_1 \cache_data_A_reg[1][8]  ( .ip(n7248), .ck(clk), .q(
        \cache_data_A[1][8] ) );
  dp_1 \cache_data_A_reg[1][9]  ( .ip(n7247), .ck(clk), .q(
        \cache_data_A[1][9] ) );
  dp_1 \cache_data_A_reg[1][10]  ( .ip(n7246), .ck(clk), .q(
        \cache_data_A[1][10] ) );
  dp_1 \cache_data_A_reg[1][11]  ( .ip(n7245), .ck(clk), .q(
        \cache_data_A[1][11] ) );
  dp_1 \cache_data_A_reg[1][12]  ( .ip(n7244), .ck(clk), .q(
        \cache_data_A[1][12] ) );
  dp_1 \cache_data_A_reg[1][13]  ( .ip(n7243), .ck(clk), .q(
        \cache_data_A[1][13] ) );
  dp_1 \cache_data_A_reg[1][14]  ( .ip(n7242), .ck(clk), .q(
        \cache_data_A[1][14] ) );
  dp_1 \cache_data_A_reg[1][15]  ( .ip(n7241), .ck(clk), .q(
        \cache_data_A[1][15] ) );
  dp_1 \cache_data_A_reg[1][16]  ( .ip(n7240), .ck(clk), .q(
        \cache_data_A[1][16] ) );
  dp_1 \cache_data_A_reg[1][17]  ( .ip(n7239), .ck(clk), .q(
        \cache_data_A[1][17] ) );
  dp_1 \cache_data_A_reg[1][18]  ( .ip(n7238), .ck(clk), .q(
        \cache_data_A[1][18] ) );
  dp_1 \cache_data_A_reg[1][19]  ( .ip(n7237), .ck(clk), .q(
        \cache_data_A[1][19] ) );
  dp_1 \cache_data_A_reg[1][20]  ( .ip(n7236), .ck(clk), .q(
        \cache_data_A[1][20] ) );
  dp_1 \cache_data_A_reg[1][21]  ( .ip(n7235), .ck(clk), .q(
        \cache_data_A[1][21] ) );
  dp_1 \cache_data_A_reg[1][22]  ( .ip(n7234), .ck(clk), .q(
        \cache_data_A[1][22] ) );
  dp_1 \cache_data_A_reg[1][23]  ( .ip(n7233), .ck(clk), .q(
        \cache_data_A[1][23] ) );
  dp_1 \cache_data_A_reg[1][24]  ( .ip(n7232), .ck(clk), .q(
        \cache_data_A[1][24] ) );
  dp_1 \cache_data_A_reg[1][25]  ( .ip(n7231), .ck(clk), .q(
        \cache_data_A[1][25] ) );
  dp_1 \cache_data_A_reg[1][26]  ( .ip(n7230), .ck(clk), .q(
        \cache_data_A[1][26] ) );
  dp_1 \cache_data_A_reg[1][27]  ( .ip(n7229), .ck(clk), .q(
        \cache_data_A[1][27] ) );
  dp_1 \cache_data_A_reg[1][28]  ( .ip(n7228), .ck(clk), .q(
        \cache_data_A[1][28] ) );
  dp_1 \cache_data_A_reg[1][29]  ( .ip(n7227), .ck(clk), .q(
        \cache_data_A[1][29] ) );
  dp_1 \cache_data_A_reg[1][30]  ( .ip(n7226), .ck(clk), .q(
        \cache_data_A[1][30] ) );
  dp_1 \cache_data_A_reg[1][31]  ( .ip(n7225), .ck(clk), .q(
        \cache_data_A[1][31] ) );
  dp_1 \cache_data_A_reg[2][0]  ( .ip(n7128), .ck(clk), .q(
        \cache_data_A[2][0] ) );
  dp_1 \cache_data_A_reg[2][1]  ( .ip(n7127), .ck(clk), .q(
        \cache_data_A[2][1] ) );
  dp_1 \cache_data_A_reg[2][2]  ( .ip(n7126), .ck(clk), .q(
        \cache_data_A[2][2] ) );
  dp_1 \cache_data_A_reg[2][3]  ( .ip(n7125), .ck(clk), .q(
        \cache_data_A[2][3] ) );
  dp_1 \cache_data_A_reg[2][4]  ( .ip(n7124), .ck(clk), .q(
        \cache_data_A[2][4] ) );
  dp_1 \cache_data_A_reg[2][5]  ( .ip(n7123), .ck(clk), .q(
        \cache_data_A[2][5] ) );
  dp_1 \cache_data_A_reg[2][6]  ( .ip(n7122), .ck(clk), .q(
        \cache_data_A[2][6] ) );
  dp_1 \cache_data_A_reg[2][7]  ( .ip(n7121), .ck(clk), .q(
        \cache_data_A[2][7] ) );
  dp_1 \cache_data_A_reg[2][8]  ( .ip(n7120), .ck(clk), .q(
        \cache_data_A[2][8] ) );
  dp_1 \cache_data_A_reg[2][9]  ( .ip(n7119), .ck(clk), .q(
        \cache_data_A[2][9] ) );
  dp_1 \cache_data_A_reg[2][10]  ( .ip(n7118), .ck(clk), .q(
        \cache_data_A[2][10] ) );
  dp_1 \cache_data_A_reg[2][11]  ( .ip(n7117), .ck(clk), .q(
        \cache_data_A[2][11] ) );
  dp_1 \cache_data_A_reg[2][12]  ( .ip(n7116), .ck(clk), .q(
        \cache_data_A[2][12] ) );
  dp_1 \cache_data_A_reg[2][13]  ( .ip(n7115), .ck(clk), .q(
        \cache_data_A[2][13] ) );
  dp_1 \cache_data_A_reg[2][14]  ( .ip(n7114), .ck(clk), .q(
        \cache_data_A[2][14] ) );
  dp_1 \cache_data_A_reg[2][15]  ( .ip(n7113), .ck(clk), .q(
        \cache_data_A[2][15] ) );
  dp_1 \cache_data_A_reg[2][16]  ( .ip(n7112), .ck(clk), .q(
        \cache_data_A[2][16] ) );
  dp_1 \cache_data_A_reg[2][17]  ( .ip(n7111), .ck(clk), .q(
        \cache_data_A[2][17] ) );
  dp_1 \cache_data_A_reg[2][18]  ( .ip(n7110), .ck(clk), .q(
        \cache_data_A[2][18] ) );
  dp_1 \cache_data_A_reg[2][19]  ( .ip(n7109), .ck(clk), .q(
        \cache_data_A[2][19] ) );
  dp_1 \cache_data_A_reg[2][20]  ( .ip(n7108), .ck(clk), .q(
        \cache_data_A[2][20] ) );
  dp_1 \cache_data_A_reg[2][21]  ( .ip(n7107), .ck(clk), .q(
        \cache_data_A[2][21] ) );
  dp_1 \cache_data_A_reg[2][22]  ( .ip(n7106), .ck(clk), .q(
        \cache_data_A[2][22] ) );
  dp_1 \cache_data_A_reg[2][23]  ( .ip(n7105), .ck(clk), .q(
        \cache_data_A[2][23] ) );
  dp_1 \cache_data_A_reg[2][24]  ( .ip(n7104), .ck(clk), .q(
        \cache_data_A[2][24] ) );
  dp_1 \cache_data_A_reg[2][25]  ( .ip(n7103), .ck(clk), .q(
        \cache_data_A[2][25] ) );
  dp_1 \cache_data_A_reg[2][26]  ( .ip(n7102), .ck(clk), .q(
        \cache_data_A[2][26] ) );
  dp_1 \cache_data_A_reg[2][27]  ( .ip(n7101), .ck(clk), .q(
        \cache_data_A[2][27] ) );
  dp_1 \cache_data_A_reg[2][28]  ( .ip(n7100), .ck(clk), .q(
        \cache_data_A[2][28] ) );
  dp_1 \cache_data_A_reg[2][29]  ( .ip(n7099), .ck(clk), .q(
        \cache_data_A[2][29] ) );
  dp_1 \cache_data_A_reg[2][30]  ( .ip(n7098), .ck(clk), .q(
        \cache_data_A[2][30] ) );
  dp_1 \cache_data_A_reg[2][31]  ( .ip(n7097), .ck(clk), .q(
        \cache_data_A[2][31] ) );
  dp_1 \cache_data_A_reg[3][0]  ( .ip(n7000), .ck(clk), .q(
        \cache_data_A[3][0] ) );
  dp_1 \cache_data_A_reg[3][1]  ( .ip(n6999), .ck(clk), .q(
        \cache_data_A[3][1] ) );
  dp_1 \cache_data_A_reg[3][2]  ( .ip(n6998), .ck(clk), .q(
        \cache_data_A[3][2] ) );
  dp_1 \cache_data_A_reg[3][3]  ( .ip(n6997), .ck(clk), .q(
        \cache_data_A[3][3] ) );
  dp_1 \cache_data_A_reg[3][4]  ( .ip(n6996), .ck(clk), .q(
        \cache_data_A[3][4] ) );
  dp_1 \cache_data_A_reg[3][5]  ( .ip(n6995), .ck(clk), .q(
        \cache_data_A[3][5] ) );
  dp_1 \cache_data_A_reg[3][6]  ( .ip(n6994), .ck(clk), .q(
        \cache_data_A[3][6] ) );
  dp_1 \cache_data_A_reg[3][7]  ( .ip(n6993), .ck(clk), .q(
        \cache_data_A[3][7] ) );
  dp_1 \cache_data_A_reg[3][8]  ( .ip(n6992), .ck(clk), .q(
        \cache_data_A[3][8] ) );
  dp_1 \cache_data_A_reg[3][9]  ( .ip(n6991), .ck(clk), .q(
        \cache_data_A[3][9] ) );
  dp_1 \cache_data_A_reg[3][10]  ( .ip(n6990), .ck(clk), .q(
        \cache_data_A[3][10] ) );
  dp_1 \cache_data_A_reg[3][11]  ( .ip(n6989), .ck(clk), .q(
        \cache_data_A[3][11] ) );
  dp_1 \cache_data_A_reg[3][12]  ( .ip(n6988), .ck(clk), .q(
        \cache_data_A[3][12] ) );
  dp_1 \cache_data_A_reg[3][13]  ( .ip(n6987), .ck(clk), .q(
        \cache_data_A[3][13] ) );
  dp_1 \cache_data_A_reg[3][14]  ( .ip(n6986), .ck(clk), .q(
        \cache_data_A[3][14] ) );
  dp_1 \cache_data_A_reg[3][15]  ( .ip(n6985), .ck(clk), .q(
        \cache_data_A[3][15] ) );
  dp_1 \cache_data_A_reg[3][16]  ( .ip(n6984), .ck(clk), .q(
        \cache_data_A[3][16] ) );
  dp_1 \cache_data_A_reg[3][17]  ( .ip(n6983), .ck(clk), .q(
        \cache_data_A[3][17] ) );
  dp_1 \cache_data_A_reg[3][18]  ( .ip(n6982), .ck(clk), .q(
        \cache_data_A[3][18] ) );
  dp_1 \cache_data_A_reg[3][19]  ( .ip(n6981), .ck(clk), .q(
        \cache_data_A[3][19] ) );
  dp_1 \cache_data_A_reg[3][20]  ( .ip(n6980), .ck(clk), .q(
        \cache_data_A[3][20] ) );
  dp_1 \cache_data_A_reg[3][21]  ( .ip(n6979), .ck(clk), .q(
        \cache_data_A[3][21] ) );
  dp_1 \cache_data_A_reg[3][22]  ( .ip(n6978), .ck(clk), .q(
        \cache_data_A[3][22] ) );
  dp_1 \cache_data_A_reg[3][23]  ( .ip(n6977), .ck(clk), .q(
        \cache_data_A[3][23] ) );
  dp_1 \cache_data_A_reg[3][24]  ( .ip(n6976), .ck(clk), .q(
        \cache_data_A[3][24] ) );
  dp_1 \cache_data_A_reg[3][25]  ( .ip(n6975), .ck(clk), .q(
        \cache_data_A[3][25] ) );
  dp_1 \cache_data_A_reg[3][26]  ( .ip(n6974), .ck(clk), .q(
        \cache_data_A[3][26] ) );
  dp_1 \cache_data_A_reg[3][27]  ( .ip(n6973), .ck(clk), .q(
        \cache_data_A[3][27] ) );
  dp_1 \cache_data_A_reg[3][28]  ( .ip(n6972), .ck(clk), .q(
        \cache_data_A[3][28] ) );
  dp_1 \cache_data_A_reg[3][29]  ( .ip(n6971), .ck(clk), .q(
        \cache_data_A[3][29] ) );
  dp_1 \cache_data_A_reg[3][30]  ( .ip(n6970), .ck(clk), .q(
        \cache_data_A[3][30] ) );
  dp_1 \cache_data_A_reg[3][31]  ( .ip(n6969), .ck(clk), .q(
        \cache_data_A[3][31] ) );
  dp_1 \cache_data_A_reg[4][8]  ( .ip(n6872), .ck(clk), .q(
        \cache_data_A[4][8] ) );
  dp_1 \cache_data_A_reg[4][9]  ( .ip(n6871), .ck(clk), .q(
        \cache_data_A[4][9] ) );
  dp_1 \cache_data_A_reg[4][10]  ( .ip(n6870), .ck(clk), .q(
        \cache_data_A[4][10] ) );
  dp_1 \cache_data_A_reg[4][11]  ( .ip(n6869), .ck(clk), .q(
        \cache_data_A[4][11] ) );
  dp_1 \cache_data_A_reg[4][12]  ( .ip(n6868), .ck(clk), .q(
        \cache_data_A[4][12] ) );
  dp_1 \cache_data_A_reg[4][13]  ( .ip(n6867), .ck(clk), .q(
        \cache_data_A[4][13] ) );
  dp_1 \cache_data_A_reg[4][14]  ( .ip(n6866), .ck(clk), .q(
        \cache_data_A[4][14] ) );
  dp_1 \cache_data_A_reg[4][15]  ( .ip(n6865), .ck(clk), .q(
        \cache_data_A[4][15] ) );
  dp_1 \cache_data_A_reg[4][16]  ( .ip(n6864), .ck(clk), .q(
        \cache_data_A[4][16] ) );
  dp_1 \cache_data_A_reg[4][17]  ( .ip(n6863), .ck(clk), .q(
        \cache_data_A[4][17] ) );
  dp_1 \cache_data_A_reg[4][18]  ( .ip(n6862), .ck(clk), .q(
        \cache_data_A[4][18] ) );
  dp_1 \cache_data_A_reg[4][19]  ( .ip(n6861), .ck(clk), .q(
        \cache_data_A[4][19] ) );
  dp_1 \cache_data_A_reg[4][20]  ( .ip(n6860), .ck(clk), .q(
        \cache_data_A[4][20] ) );
  dp_1 \cache_data_A_reg[4][21]  ( .ip(n6859), .ck(clk), .q(
        \cache_data_A[4][21] ) );
  dp_1 \cache_data_A_reg[4][22]  ( .ip(n6858), .ck(clk), .q(
        \cache_data_A[4][22] ) );
  dp_1 \cache_data_A_reg[4][23]  ( .ip(n6857), .ck(clk), .q(
        \cache_data_A[4][23] ) );
  dp_1 \cache_data_A_reg[4][24]  ( .ip(n6856), .ck(clk), .q(
        \cache_data_A[4][24] ) );
  dp_1 \cache_data_A_reg[4][25]  ( .ip(n6855), .ck(clk), .q(
        \cache_data_A[4][25] ) );
  dp_1 \cache_data_A_reg[4][26]  ( .ip(n6854), .ck(clk), .q(
        \cache_data_A[4][26] ) );
  dp_1 \cache_data_A_reg[4][27]  ( .ip(n6853), .ck(clk), .q(
        \cache_data_A[4][27] ) );
  dp_1 \cache_data_A_reg[4][28]  ( .ip(n6852), .ck(clk), .q(
        \cache_data_A[4][28] ) );
  dp_1 \cache_data_A_reg[4][29]  ( .ip(n6851), .ck(clk), .q(
        \cache_data_A[4][29] ) );
  dp_1 \cache_data_A_reg[4][30]  ( .ip(n6850), .ck(clk), .q(
        \cache_data_A[4][30] ) );
  dp_1 \cache_data_A_reg[4][31]  ( .ip(n6849), .ck(clk), .q(
        \cache_data_A[4][31] ) );
  dp_1 \cache_data_A_reg[4][0]  ( .ip(n6848), .ck(clk), .q(
        \cache_data_A[4][0] ) );
  dp_1 \cache_data_A_reg[4][1]  ( .ip(n6847), .ck(clk), .q(
        \cache_data_A[4][1] ) );
  dp_1 \cache_data_A_reg[4][2]  ( .ip(n6846), .ck(clk), .q(
        \cache_data_A[4][2] ) );
  dp_1 \cache_data_A_reg[4][3]  ( .ip(n6845), .ck(clk), .q(
        \cache_data_A[4][3] ) );
  dp_1 \cache_data_A_reg[4][4]  ( .ip(n6844), .ck(clk), .q(
        \cache_data_A[4][4] ) );
  dp_1 \cache_data_A_reg[4][5]  ( .ip(n6843), .ck(clk), .q(
        \cache_data_A[4][5] ) );
  dp_1 \cache_data_A_reg[4][6]  ( .ip(n6842), .ck(clk), .q(
        \cache_data_A[4][6] ) );
  dp_1 \cache_data_A_reg[4][7]  ( .ip(n6841), .ck(clk), .q(
        \cache_data_A[4][7] ) );
  dp_1 \cache_data_A_reg[5][0]  ( .ip(n6744), .ck(clk), .q(
        \cache_data_A[5][0] ) );
  dp_1 \cache_data_A_reg[5][1]  ( .ip(n6743), .ck(clk), .q(
        \cache_data_A[5][1] ) );
  dp_1 \cache_data_A_reg[5][2]  ( .ip(n6742), .ck(clk), .q(
        \cache_data_A[5][2] ) );
  dp_1 \cache_data_A_reg[5][3]  ( .ip(n6741), .ck(clk), .q(
        \cache_data_A[5][3] ) );
  dp_1 \cache_data_A_reg[5][4]  ( .ip(n6740), .ck(clk), .q(
        \cache_data_A[5][4] ) );
  dp_1 \cache_data_A_reg[5][5]  ( .ip(n6739), .ck(clk), .q(
        \cache_data_A[5][5] ) );
  dp_1 \cache_data_A_reg[5][6]  ( .ip(n6738), .ck(clk), .q(
        \cache_data_A[5][6] ) );
  dp_1 \cache_data_A_reg[5][7]  ( .ip(n6737), .ck(clk), .q(
        \cache_data_A[5][7] ) );
  dp_1 \cache_data_A_reg[5][8]  ( .ip(n6736), .ck(clk), .q(
        \cache_data_A[5][8] ) );
  dp_1 \cache_data_A_reg[5][9]  ( .ip(n6735), .ck(clk), .q(
        \cache_data_A[5][9] ) );
  dp_1 \cache_data_A_reg[5][10]  ( .ip(n6734), .ck(clk), .q(
        \cache_data_A[5][10] ) );
  dp_1 \cache_data_A_reg[5][11]  ( .ip(n6733), .ck(clk), .q(
        \cache_data_A[5][11] ) );
  dp_1 \cache_data_A_reg[5][12]  ( .ip(n6732), .ck(clk), .q(
        \cache_data_A[5][12] ) );
  dp_1 \cache_data_A_reg[5][13]  ( .ip(n6731), .ck(clk), .q(
        \cache_data_A[5][13] ) );
  dp_1 \cache_data_A_reg[5][14]  ( .ip(n6730), .ck(clk), .q(
        \cache_data_A[5][14] ) );
  dp_1 \cache_data_A_reg[5][15]  ( .ip(n6729), .ck(clk), .q(
        \cache_data_A[5][15] ) );
  dp_1 \cache_data_A_reg[5][16]  ( .ip(n6728), .ck(clk), .q(
        \cache_data_A[5][16] ) );
  dp_1 \cache_data_A_reg[5][17]  ( .ip(n6727), .ck(clk), .q(
        \cache_data_A[5][17] ) );
  dp_1 \cache_data_A_reg[5][18]  ( .ip(n6726), .ck(clk), .q(
        \cache_data_A[5][18] ) );
  dp_1 \cache_data_A_reg[5][19]  ( .ip(n6725), .ck(clk), .q(
        \cache_data_A[5][19] ) );
  dp_1 \cache_data_A_reg[5][20]  ( .ip(n6724), .ck(clk), .q(
        \cache_data_A[5][20] ) );
  dp_1 \cache_data_A_reg[5][21]  ( .ip(n6723), .ck(clk), .q(
        \cache_data_A[5][21] ) );
  dp_1 \cache_data_A_reg[5][22]  ( .ip(n6722), .ck(clk), .q(
        \cache_data_A[5][22] ) );
  dp_1 \cache_data_A_reg[5][23]  ( .ip(n6721), .ck(clk), .q(
        \cache_data_A[5][23] ) );
  dp_1 \cache_data_A_reg[5][24]  ( .ip(n6720), .ck(clk), .q(
        \cache_data_A[5][24] ) );
  dp_1 \cache_data_A_reg[5][25]  ( .ip(n6719), .ck(clk), .q(
        \cache_data_A[5][25] ) );
  dp_1 \cache_data_A_reg[5][26]  ( .ip(n6718), .ck(clk), .q(
        \cache_data_A[5][26] ) );
  dp_1 \cache_data_A_reg[5][27]  ( .ip(n6717), .ck(clk), .q(
        \cache_data_A[5][27] ) );
  dp_1 \cache_data_A_reg[5][28]  ( .ip(n6716), .ck(clk), .q(
        \cache_data_A[5][28] ) );
  dp_1 \cache_data_A_reg[5][29]  ( .ip(n6715), .ck(clk), .q(
        \cache_data_A[5][29] ) );
  dp_1 \cache_data_A_reg[5][30]  ( .ip(n6714), .ck(clk), .q(
        \cache_data_A[5][30] ) );
  dp_1 \cache_data_A_reg[5][31]  ( .ip(n6713), .ck(clk), .q(
        \cache_data_A[5][31] ) );
  dp_1 \cache_data_A_reg[6][0]  ( .ip(n6616), .ck(clk), .q(
        \cache_data_A[6][0] ) );
  dp_1 \cache_data_A_reg[6][1]  ( .ip(n6615), .ck(clk), .q(
        \cache_data_A[6][1] ) );
  dp_1 \cache_data_A_reg[6][2]  ( .ip(n6614), .ck(clk), .q(
        \cache_data_A[6][2] ) );
  dp_1 \cache_data_A_reg[6][3]  ( .ip(n6613), .ck(clk), .q(
        \cache_data_A[6][3] ) );
  dp_1 \cache_data_A_reg[6][4]  ( .ip(n6612), .ck(clk), .q(
        \cache_data_A[6][4] ) );
  dp_1 \cache_data_A_reg[6][5]  ( .ip(n6611), .ck(clk), .q(
        \cache_data_A[6][5] ) );
  dp_1 \cache_data_A_reg[6][6]  ( .ip(n6610), .ck(clk), .q(
        \cache_data_A[6][6] ) );
  dp_1 \cache_data_A_reg[6][7]  ( .ip(n6609), .ck(clk), .q(
        \cache_data_A[6][7] ) );
  dp_1 \cache_data_A_reg[6][8]  ( .ip(n6608), .ck(clk), .q(
        \cache_data_A[6][8] ) );
  dp_1 \cache_data_A_reg[6][9]  ( .ip(n6607), .ck(clk), .q(
        \cache_data_A[6][9] ) );
  dp_1 \cache_data_A_reg[6][10]  ( .ip(n6606), .ck(clk), .q(
        \cache_data_A[6][10] ) );
  dp_1 \cache_data_A_reg[6][11]  ( .ip(n6605), .ck(clk), .q(
        \cache_data_A[6][11] ) );
  dp_1 \cache_data_A_reg[6][12]  ( .ip(n6604), .ck(clk), .q(
        \cache_data_A[6][12] ) );
  dp_1 \cache_data_A_reg[6][13]  ( .ip(n6603), .ck(clk), .q(
        \cache_data_A[6][13] ) );
  dp_1 \cache_data_A_reg[6][14]  ( .ip(n6602), .ck(clk), .q(
        \cache_data_A[6][14] ) );
  dp_1 \cache_data_A_reg[6][15]  ( .ip(n6601), .ck(clk), .q(
        \cache_data_A[6][15] ) );
  dp_1 \cache_data_A_reg[6][16]  ( .ip(n6600), .ck(clk), .q(
        \cache_data_A[6][16] ) );
  dp_1 \cache_data_A_reg[6][17]  ( .ip(n6599), .ck(clk), .q(
        \cache_data_A[6][17] ) );
  dp_1 \cache_data_A_reg[6][18]  ( .ip(n6598), .ck(clk), .q(
        \cache_data_A[6][18] ) );
  dp_1 \cache_data_A_reg[6][19]  ( .ip(n6597), .ck(clk), .q(
        \cache_data_A[6][19] ) );
  dp_1 \cache_data_A_reg[6][20]  ( .ip(n6596), .ck(clk), .q(
        \cache_data_A[6][20] ) );
  dp_1 \cache_data_A_reg[6][21]  ( .ip(n6595), .ck(clk), .q(
        \cache_data_A[6][21] ) );
  dp_1 \cache_data_A_reg[6][22]  ( .ip(n6594), .ck(clk), .q(
        \cache_data_A[6][22] ) );
  dp_1 \cache_data_A_reg[6][23]  ( .ip(n6593), .ck(clk), .q(
        \cache_data_A[6][23] ) );
  dp_1 \cache_data_A_reg[6][24]  ( .ip(n6592), .ck(clk), .q(
        \cache_data_A[6][24] ) );
  dp_1 \cache_data_A_reg[6][25]  ( .ip(n6591), .ck(clk), .q(
        \cache_data_A[6][25] ) );
  dp_1 \cache_data_A_reg[6][26]  ( .ip(n6590), .ck(clk), .q(
        \cache_data_A[6][26] ) );
  dp_1 \cache_data_A_reg[6][27]  ( .ip(n6589), .ck(clk), .q(
        \cache_data_A[6][27] ) );
  dp_1 \cache_data_A_reg[6][28]  ( .ip(n6588), .ck(clk), .q(
        \cache_data_A[6][28] ) );
  dp_1 \cache_data_A_reg[6][29]  ( .ip(n6587), .ck(clk), .q(
        \cache_data_A[6][29] ) );
  dp_1 \cache_data_A_reg[6][30]  ( .ip(n6586), .ck(clk), .q(
        \cache_data_A[6][30] ) );
  dp_1 \cache_data_A_reg[6][31]  ( .ip(n6585), .ck(clk), .q(
        \cache_data_A[6][31] ) );
  dp_1 \cache_data_A_reg[7][20]  ( .ip(n6488), .ck(clk), .q(
        \cache_data_A[7][20] ) );
  dp_1 \cache_data_A_reg[7][21]  ( .ip(n6487), .ck(clk), .q(
        \cache_data_A[7][21] ) );
  dp_1 \cache_data_A_reg[7][22]  ( .ip(n6486), .ck(clk), .q(
        \cache_data_A[7][22] ) );
  dp_1 \cache_data_A_reg[7][23]  ( .ip(n6485), .ck(clk), .q(
        \cache_data_A[7][23] ) );
  dp_1 \cache_data_A_reg[7][24]  ( .ip(n6484), .ck(clk), .q(
        \cache_data_A[7][24] ) );
  dp_1 \cache_data_A_reg[7][25]  ( .ip(n6483), .ck(clk), .q(
        \cache_data_A[7][25] ) );
  dp_1 \cache_data_A_reg[7][26]  ( .ip(n6482), .ck(clk), .q(
        \cache_data_A[7][26] ) );
  dp_1 \cache_data_A_reg[7][27]  ( .ip(n6481), .ck(clk), .q(
        \cache_data_A[7][27] ) );
  dp_1 \cache_data_A_reg[7][28]  ( .ip(n6480), .ck(clk), .q(
        \cache_data_A[7][28] ) );
  dp_1 \cache_data_A_reg[7][29]  ( .ip(n6479), .ck(clk), .q(
        \cache_data_A[7][29] ) );
  dp_1 \cache_data_A_reg[7][30]  ( .ip(n6478), .ck(clk), .q(
        \cache_data_A[7][30] ) );
  dp_1 \cache_data_A_reg[7][31]  ( .ip(n6477), .ck(clk), .q(
        \cache_data_A[7][31] ) );
  dp_1 \cache_data_A_reg[7][0]  ( .ip(n6476), .ck(clk), .q(
        \cache_data_A[7][0] ) );
  dp_1 \cache_data_A_reg[7][1]  ( .ip(n6475), .ck(clk), .q(
        \cache_data_A[7][1] ) );
  dp_1 \cache_data_A_reg[7][2]  ( .ip(n6474), .ck(clk), .q(
        \cache_data_A[7][2] ) );
  dp_1 \cache_data_A_reg[7][3]  ( .ip(n6473), .ck(clk), .q(
        \cache_data_A[7][3] ) );
  dp_1 \cache_data_A_reg[7][4]  ( .ip(n6472), .ck(clk), .q(
        \cache_data_A[7][4] ) );
  dp_1 \cache_data_A_reg[7][5]  ( .ip(n6471), .ck(clk), .q(
        \cache_data_A[7][5] ) );
  dp_1 \cache_data_A_reg[7][6]  ( .ip(n6470), .ck(clk), .q(
        \cache_data_A[7][6] ) );
  dp_1 \cache_data_A_reg[7][7]  ( .ip(n6469), .ck(clk), .q(
        \cache_data_A[7][7] ) );
  dp_1 \cache_data_A_reg[7][8]  ( .ip(n6468), .ck(clk), .q(
        \cache_data_A[7][8] ) );
  dp_1 \cache_data_A_reg[7][9]  ( .ip(n6467), .ck(clk), .q(
        \cache_data_A[7][9] ) );
  dp_1 \cache_data_A_reg[7][10]  ( .ip(n6466), .ck(clk), .q(
        \cache_data_A[7][10] ) );
  dp_1 \cache_data_A_reg[7][11]  ( .ip(n6465), .ck(clk), .q(
        \cache_data_A[7][11] ) );
  dp_1 \cache_data_A_reg[7][12]  ( .ip(n6464), .ck(clk), .q(
        \cache_data_A[7][12] ) );
  dp_1 \cache_data_A_reg[7][13]  ( .ip(n6463), .ck(clk), .q(
        \cache_data_A[7][13] ) );
  dp_1 \cache_data_A_reg[7][14]  ( .ip(n6462), .ck(clk), .q(
        \cache_data_A[7][14] ) );
  dp_1 \cache_data_A_reg[7][15]  ( .ip(n6461), .ck(clk), .q(
        \cache_data_A[7][15] ) );
  dp_1 \cache_data_A_reg[7][16]  ( .ip(n6460), .ck(clk), .q(
        \cache_data_A[7][16] ) );
  dp_1 \cache_data_A_reg[7][17]  ( .ip(n6459), .ck(clk), .q(
        \cache_data_A[7][17] ) );
  dp_1 \cache_data_A_reg[7][18]  ( .ip(n6458), .ck(clk), .q(
        \cache_data_A[7][18] ) );
  dp_1 \cache_data_A_reg[7][19]  ( .ip(n6457), .ck(clk), .q(
        \cache_data_A[7][19] ) );
  dp_1 \cache_data_A_reg[0][32]  ( .ip(n7352), .ck(clk), .q(
        \cache_data_A[0][32] ) );
  dp_1 \cache_data_A_reg[0][33]  ( .ip(n7351), .ck(clk), .q(
        \cache_data_A[0][33] ) );
  dp_1 \cache_data_A_reg[0][34]  ( .ip(n7350), .ck(clk), .q(
        \cache_data_A[0][34] ) );
  dp_1 \cache_data_A_reg[0][35]  ( .ip(n7349), .ck(clk), .q(
        \cache_data_A[0][35] ) );
  dp_1 \cache_data_A_reg[0][36]  ( .ip(n7348), .ck(clk), .q(
        \cache_data_A[0][36] ) );
  dp_1 \cache_data_A_reg[0][37]  ( .ip(n7347), .ck(clk), .q(
        \cache_data_A[0][37] ) );
  dp_1 \cache_data_A_reg[0][38]  ( .ip(n7346), .ck(clk), .q(
        \cache_data_A[0][38] ) );
  dp_1 \cache_data_A_reg[0][39]  ( .ip(n7345), .ck(clk), .q(
        \cache_data_A[0][39] ) );
  dp_1 \cache_data_A_reg[0][40]  ( .ip(n7344), .ck(clk), .q(
        \cache_data_A[0][40] ) );
  dp_1 \cache_data_A_reg[0][41]  ( .ip(n7343), .ck(clk), .q(
        \cache_data_A[0][41] ) );
  dp_1 \cache_data_A_reg[0][42]  ( .ip(n7342), .ck(clk), .q(
        \cache_data_A[0][42] ) );
  dp_1 \cache_data_A_reg[0][43]  ( .ip(n7341), .ck(clk), .q(
        \cache_data_A[0][43] ) );
  dp_1 \cache_data_A_reg[0][44]  ( .ip(n7340), .ck(clk), .q(
        \cache_data_A[0][44] ) );
  dp_1 \cache_data_A_reg[0][45]  ( .ip(n7339), .ck(clk), .q(
        \cache_data_A[0][45] ) );
  dp_1 \cache_data_A_reg[0][46]  ( .ip(n7338), .ck(clk), .q(
        \cache_data_A[0][46] ) );
  dp_1 \cache_data_A_reg[0][47]  ( .ip(n7337), .ck(clk), .q(
        \cache_data_A[0][47] ) );
  dp_1 \cache_data_A_reg[0][48]  ( .ip(n7336), .ck(clk), .q(
        \cache_data_A[0][48] ) );
  dp_1 \cache_data_A_reg[0][49]  ( .ip(n7335), .ck(clk), .q(
        \cache_data_A[0][49] ) );
  dp_1 \cache_data_A_reg[0][50]  ( .ip(n7334), .ck(clk), .q(
        \cache_data_A[0][50] ) );
  dp_1 \cache_data_A_reg[0][51]  ( .ip(n7333), .ck(clk), .q(
        \cache_data_A[0][51] ) );
  dp_1 \cache_data_A_reg[0][52]  ( .ip(n7332), .ck(clk), .q(
        \cache_data_A[0][52] ) );
  dp_1 \cache_data_A_reg[0][53]  ( .ip(n7331), .ck(clk), .q(
        \cache_data_A[0][53] ) );
  dp_1 \cache_data_A_reg[0][54]  ( .ip(n7330), .ck(clk), .q(
        \cache_data_A[0][54] ) );
  dp_1 \cache_data_A_reg[0][55]  ( .ip(n7329), .ck(clk), .q(
        \cache_data_A[0][55] ) );
  dp_1 \cache_data_A_reg[0][56]  ( .ip(n7328), .ck(clk), .q(
        \cache_data_A[0][56] ) );
  dp_1 \cache_data_A_reg[0][57]  ( .ip(n7327), .ck(clk), .q(
        \cache_data_A[0][57] ) );
  dp_1 \cache_data_A_reg[0][58]  ( .ip(n7326), .ck(clk), .q(
        \cache_data_A[0][58] ) );
  dp_1 \cache_data_A_reg[0][59]  ( .ip(n7325), .ck(clk), .q(
        \cache_data_A[0][59] ) );
  dp_1 \cache_data_A_reg[0][60]  ( .ip(n7324), .ck(clk), .q(
        \cache_data_A[0][60] ) );
  dp_1 \cache_data_A_reg[0][61]  ( .ip(n7323), .ck(clk), .q(
        \cache_data_A[0][61] ) );
  dp_1 \cache_data_A_reg[0][62]  ( .ip(n7322), .ck(clk), .q(
        \cache_data_A[0][62] ) );
  dp_1 \cache_data_A_reg[0][63]  ( .ip(n7321), .ck(clk), .q(
        \cache_data_A[0][63] ) );
  dp_1 \cache_data_A_reg[1][32]  ( .ip(n7224), .ck(clk), .q(
        \cache_data_A[1][32] ) );
  dp_1 \cache_data_A_reg[1][33]  ( .ip(n7223), .ck(clk), .q(
        \cache_data_A[1][33] ) );
  dp_1 \cache_data_A_reg[1][34]  ( .ip(n7222), .ck(clk), .q(
        \cache_data_A[1][34] ) );
  dp_1 \cache_data_A_reg[1][35]  ( .ip(n7221), .ck(clk), .q(
        \cache_data_A[1][35] ) );
  dp_1 \cache_data_A_reg[1][36]  ( .ip(n7220), .ck(clk), .q(
        \cache_data_A[1][36] ) );
  dp_1 \cache_data_A_reg[1][37]  ( .ip(n7219), .ck(clk), .q(
        \cache_data_A[1][37] ) );
  dp_1 \cache_data_A_reg[1][38]  ( .ip(n7218), .ck(clk), .q(
        \cache_data_A[1][38] ) );
  dp_1 \cache_data_A_reg[1][39]  ( .ip(n7217), .ck(clk), .q(
        \cache_data_A[1][39] ) );
  dp_1 \cache_data_A_reg[1][40]  ( .ip(n7216), .ck(clk), .q(
        \cache_data_A[1][40] ) );
  dp_1 \cache_data_A_reg[1][41]  ( .ip(n7215), .ck(clk), .q(
        \cache_data_A[1][41] ) );
  dp_1 \cache_data_A_reg[1][42]  ( .ip(n7214), .ck(clk), .q(
        \cache_data_A[1][42] ) );
  dp_1 \cache_data_A_reg[1][43]  ( .ip(n7213), .ck(clk), .q(
        \cache_data_A[1][43] ) );
  dp_1 \cache_data_A_reg[1][44]  ( .ip(n7212), .ck(clk), .q(
        \cache_data_A[1][44] ) );
  dp_1 \cache_data_A_reg[1][45]  ( .ip(n7211), .ck(clk), .q(
        \cache_data_A[1][45] ) );
  dp_1 \cache_data_A_reg[1][46]  ( .ip(n7210), .ck(clk), .q(
        \cache_data_A[1][46] ) );
  dp_1 \cache_data_A_reg[1][47]  ( .ip(n7209), .ck(clk), .q(
        \cache_data_A[1][47] ) );
  dp_1 \cache_data_A_reg[1][48]  ( .ip(n7208), .ck(clk), .q(
        \cache_data_A[1][48] ) );
  dp_1 \cache_data_A_reg[1][49]  ( .ip(n7207), .ck(clk), .q(
        \cache_data_A[1][49] ) );
  dp_1 \cache_data_A_reg[1][50]  ( .ip(n7206), .ck(clk), .q(
        \cache_data_A[1][50] ) );
  dp_1 \cache_data_A_reg[1][51]  ( .ip(n7205), .ck(clk), .q(
        \cache_data_A[1][51] ) );
  dp_1 \cache_data_A_reg[1][52]  ( .ip(n7204), .ck(clk), .q(
        \cache_data_A[1][52] ) );
  dp_1 \cache_data_A_reg[1][53]  ( .ip(n7203), .ck(clk), .q(
        \cache_data_A[1][53] ) );
  dp_1 \cache_data_A_reg[1][54]  ( .ip(n7202), .ck(clk), .q(
        \cache_data_A[1][54] ) );
  dp_1 \cache_data_A_reg[1][55]  ( .ip(n7201), .ck(clk), .q(
        \cache_data_A[1][55] ) );
  dp_1 \cache_data_A_reg[1][56]  ( .ip(n7200), .ck(clk), .q(
        \cache_data_A[1][56] ) );
  dp_1 \cache_data_A_reg[1][57]  ( .ip(n7199), .ck(clk), .q(
        \cache_data_A[1][57] ) );
  dp_1 \cache_data_A_reg[1][58]  ( .ip(n7198), .ck(clk), .q(
        \cache_data_A[1][58] ) );
  dp_1 \cache_data_A_reg[1][59]  ( .ip(n7197), .ck(clk), .q(
        \cache_data_A[1][59] ) );
  dp_1 \cache_data_A_reg[1][60]  ( .ip(n7196), .ck(clk), .q(
        \cache_data_A[1][60] ) );
  dp_1 \cache_data_A_reg[1][61]  ( .ip(n7195), .ck(clk), .q(
        \cache_data_A[1][61] ) );
  dp_1 \cache_data_A_reg[1][62]  ( .ip(n7194), .ck(clk), .q(
        \cache_data_A[1][62] ) );
  dp_1 \cache_data_A_reg[1][63]  ( .ip(n7193), .ck(clk), .q(
        \cache_data_A[1][63] ) );
  dp_1 \cache_data_A_reg[2][32]  ( .ip(n7096), .ck(clk), .q(
        \cache_data_A[2][32] ) );
  dp_1 \cache_data_A_reg[2][33]  ( .ip(n7095), .ck(clk), .q(
        \cache_data_A[2][33] ) );
  dp_1 \cache_data_A_reg[2][34]  ( .ip(n7094), .ck(clk), .q(
        \cache_data_A[2][34] ) );
  dp_1 \cache_data_A_reg[2][35]  ( .ip(n7093), .ck(clk), .q(
        \cache_data_A[2][35] ) );
  dp_1 \cache_data_A_reg[2][36]  ( .ip(n7092), .ck(clk), .q(
        \cache_data_A[2][36] ) );
  dp_1 \cache_data_A_reg[2][37]  ( .ip(n7091), .ck(clk), .q(
        \cache_data_A[2][37] ) );
  dp_1 \cache_data_A_reg[2][38]  ( .ip(n7090), .ck(clk), .q(
        \cache_data_A[2][38] ) );
  dp_1 \cache_data_A_reg[2][39]  ( .ip(n7089), .ck(clk), .q(
        \cache_data_A[2][39] ) );
  dp_1 \cache_data_A_reg[2][40]  ( .ip(n7088), .ck(clk), .q(
        \cache_data_A[2][40] ) );
  dp_1 \cache_data_A_reg[2][41]  ( .ip(n7087), .ck(clk), .q(
        \cache_data_A[2][41] ) );
  dp_1 \cache_data_A_reg[2][42]  ( .ip(n7086), .ck(clk), .q(
        \cache_data_A[2][42] ) );
  dp_1 \cache_data_A_reg[2][43]  ( .ip(n7085), .ck(clk), .q(
        \cache_data_A[2][43] ) );
  dp_1 \cache_data_A_reg[2][44]  ( .ip(n7084), .ck(clk), .q(
        \cache_data_A[2][44] ) );
  dp_1 \cache_data_A_reg[2][45]  ( .ip(n7083), .ck(clk), .q(
        \cache_data_A[2][45] ) );
  dp_1 \cache_data_A_reg[2][46]  ( .ip(n7082), .ck(clk), .q(
        \cache_data_A[2][46] ) );
  dp_1 \cache_data_A_reg[2][47]  ( .ip(n7081), .ck(clk), .q(
        \cache_data_A[2][47] ) );
  dp_1 \cache_data_A_reg[2][48]  ( .ip(n7080), .ck(clk), .q(
        \cache_data_A[2][48] ) );
  dp_1 \cache_data_A_reg[2][49]  ( .ip(n7079), .ck(clk), .q(
        \cache_data_A[2][49] ) );
  dp_1 \cache_data_A_reg[2][50]  ( .ip(n7078), .ck(clk), .q(
        \cache_data_A[2][50] ) );
  dp_1 \cache_data_A_reg[2][51]  ( .ip(n7077), .ck(clk), .q(
        \cache_data_A[2][51] ) );
  dp_1 \cache_data_A_reg[2][52]  ( .ip(n7076), .ck(clk), .q(
        \cache_data_A[2][52] ) );
  dp_1 \cache_data_A_reg[2][53]  ( .ip(n7075), .ck(clk), .q(
        \cache_data_A[2][53] ) );
  dp_1 \cache_data_A_reg[2][54]  ( .ip(n7074), .ck(clk), .q(
        \cache_data_A[2][54] ) );
  dp_1 \cache_data_A_reg[2][55]  ( .ip(n7073), .ck(clk), .q(
        \cache_data_A[2][55] ) );
  dp_1 \cache_data_A_reg[2][56]  ( .ip(n7072), .ck(clk), .q(
        \cache_data_A[2][56] ) );
  dp_1 \cache_data_A_reg[2][57]  ( .ip(n7071), .ck(clk), .q(
        \cache_data_A[2][57] ) );
  dp_1 \cache_data_A_reg[2][58]  ( .ip(n7070), .ck(clk), .q(
        \cache_data_A[2][58] ) );
  dp_1 \cache_data_A_reg[2][59]  ( .ip(n7069), .ck(clk), .q(
        \cache_data_A[2][59] ) );
  dp_1 \cache_data_A_reg[2][60]  ( .ip(n7068), .ck(clk), .q(
        \cache_data_A[2][60] ) );
  dp_1 \cache_data_A_reg[2][61]  ( .ip(n7067), .ck(clk), .q(
        \cache_data_A[2][61] ) );
  dp_1 \cache_data_A_reg[2][62]  ( .ip(n7066), .ck(clk), .q(
        \cache_data_A[2][62] ) );
  dp_1 \cache_data_A_reg[2][63]  ( .ip(n7065), .ck(clk), .q(
        \cache_data_A[2][63] ) );
  dp_1 \cache_data_A_reg[3][37]  ( .ip(n6968), .ck(clk), .q(
        \cache_data_A[3][37] ) );
  dp_1 \cache_data_A_reg[3][38]  ( .ip(n6967), .ck(clk), .q(
        \cache_data_A[3][38] ) );
  dp_1 \cache_data_A_reg[3][39]  ( .ip(n6966), .ck(clk), .q(
        \cache_data_A[3][39] ) );
  dp_1 \cache_data_A_reg[3][40]  ( .ip(n6965), .ck(clk), .q(
        \cache_data_A[3][40] ) );
  dp_1 \cache_data_A_reg[3][41]  ( .ip(n6964), .ck(clk), .q(
        \cache_data_A[3][41] ) );
  dp_1 \cache_data_A_reg[3][42]  ( .ip(n6963), .ck(clk), .q(
        \cache_data_A[3][42] ) );
  dp_1 \cache_data_A_reg[3][43]  ( .ip(n6962), .ck(clk), .q(
        \cache_data_A[3][43] ) );
  dp_1 \cache_data_A_reg[3][44]  ( .ip(n6961), .ck(clk), .q(
        \cache_data_A[3][44] ) );
  dp_1 \cache_data_A_reg[3][45]  ( .ip(n6960), .ck(clk), .q(
        \cache_data_A[3][45] ) );
  dp_1 \cache_data_A_reg[3][46]  ( .ip(n6959), .ck(clk), .q(
        \cache_data_A[3][46] ) );
  dp_1 \cache_data_A_reg[3][47]  ( .ip(n6958), .ck(clk), .q(
        \cache_data_A[3][47] ) );
  dp_1 \cache_data_A_reg[3][48]  ( .ip(n6957), .ck(clk), .q(
        \cache_data_A[3][48] ) );
  dp_1 \cache_data_A_reg[3][49]  ( .ip(n6956), .ck(clk), .q(
        \cache_data_A[3][49] ) );
  dp_1 \cache_data_A_reg[3][50]  ( .ip(n6955), .ck(clk), .q(
        \cache_data_A[3][50] ) );
  dp_1 \cache_data_A_reg[3][51]  ( .ip(n6954), .ck(clk), .q(
        \cache_data_A[3][51] ) );
  dp_1 \cache_data_A_reg[3][52]  ( .ip(n6953), .ck(clk), .q(
        \cache_data_A[3][52] ) );
  dp_1 \cache_data_A_reg[3][53]  ( .ip(n6952), .ck(clk), .q(
        \cache_data_A[3][53] ) );
  dp_1 \cache_data_A_reg[3][54]  ( .ip(n6951), .ck(clk), .q(
        \cache_data_A[3][54] ) );
  dp_1 \cache_data_A_reg[3][55]  ( .ip(n6950), .ck(clk), .q(
        \cache_data_A[3][55] ) );
  dp_1 \cache_data_A_reg[3][56]  ( .ip(n6949), .ck(clk), .q(
        \cache_data_A[3][56] ) );
  dp_1 \cache_data_A_reg[3][57]  ( .ip(n6948), .ck(clk), .q(
        \cache_data_A[3][57] ) );
  dp_1 \cache_data_A_reg[3][58]  ( .ip(n6947), .ck(clk), .q(
        \cache_data_A[3][58] ) );
  dp_1 \cache_data_A_reg[3][59]  ( .ip(n6946), .ck(clk), .q(
        \cache_data_A[3][59] ) );
  dp_1 \cache_data_A_reg[3][60]  ( .ip(n6945), .ck(clk), .q(
        \cache_data_A[3][60] ) );
  dp_1 \cache_data_A_reg[3][61]  ( .ip(n6944), .ck(clk), .q(
        \cache_data_A[3][61] ) );
  dp_1 \cache_data_A_reg[3][62]  ( .ip(n6943), .ck(clk), .q(
        \cache_data_A[3][62] ) );
  dp_1 \cache_data_A_reg[3][63]  ( .ip(n6942), .ck(clk), .q(
        \cache_data_A[3][63] ) );
  dp_1 \cache_data_A_reg[3][32]  ( .ip(n6941), .ck(clk), .q(
        \cache_data_A[3][32] ) );
  dp_1 \cache_data_A_reg[3][33]  ( .ip(n6940), .ck(clk), .q(
        \cache_data_A[3][33] ) );
  dp_1 \cache_data_A_reg[3][34]  ( .ip(n6939), .ck(clk), .q(
        \cache_data_A[3][34] ) );
  dp_1 \cache_data_A_reg[3][35]  ( .ip(n6938), .ck(clk), .q(
        \cache_data_A[3][35] ) );
  dp_1 \cache_data_A_reg[3][36]  ( .ip(n6937), .ck(clk), .q(
        \cache_data_A[3][36] ) );
  dp_1 \cache_data_A_reg[4][32]  ( .ip(n6840), .ck(clk), .q(
        \cache_data_A[4][32] ) );
  dp_1 \cache_data_A_reg[4][33]  ( .ip(n6839), .ck(clk), .q(
        \cache_data_A[4][33] ) );
  dp_1 \cache_data_A_reg[4][34]  ( .ip(n6838), .ck(clk), .q(
        \cache_data_A[4][34] ) );
  dp_1 \cache_data_A_reg[4][35]  ( .ip(n6837), .ck(clk), .q(
        \cache_data_A[4][35] ) );
  dp_1 \cache_data_A_reg[4][36]  ( .ip(n6836), .ck(clk), .q(
        \cache_data_A[4][36] ) );
  dp_1 \cache_data_A_reg[4][37]  ( .ip(n6835), .ck(clk), .q(
        \cache_data_A[4][37] ) );
  dp_1 \cache_data_A_reg[4][38]  ( .ip(n6834), .ck(clk), .q(
        \cache_data_A[4][38] ) );
  dp_1 \cache_data_A_reg[4][39]  ( .ip(n6833), .ck(clk), .q(
        \cache_data_A[4][39] ) );
  dp_1 \cache_data_A_reg[4][40]  ( .ip(n6832), .ck(clk), .q(
        \cache_data_A[4][40] ) );
  dp_1 \cache_data_A_reg[4][41]  ( .ip(n6831), .ck(clk), .q(
        \cache_data_A[4][41] ) );
  dp_1 \cache_data_A_reg[4][42]  ( .ip(n6830), .ck(clk), .q(
        \cache_data_A[4][42] ) );
  dp_1 \cache_data_A_reg[4][43]  ( .ip(n6829), .ck(clk), .q(
        \cache_data_A[4][43] ) );
  dp_1 \cache_data_A_reg[4][44]  ( .ip(n6828), .ck(clk), .q(
        \cache_data_A[4][44] ) );
  dp_1 \cache_data_A_reg[4][45]  ( .ip(n6827), .ck(clk), .q(
        \cache_data_A[4][45] ) );
  dp_1 \cache_data_A_reg[4][46]  ( .ip(n6826), .ck(clk), .q(
        \cache_data_A[4][46] ) );
  dp_1 \cache_data_A_reg[4][47]  ( .ip(n6825), .ck(clk), .q(
        \cache_data_A[4][47] ) );
  dp_1 \cache_data_A_reg[4][48]  ( .ip(n6824), .ck(clk), .q(
        \cache_data_A[4][48] ) );
  dp_1 \cache_data_A_reg[4][49]  ( .ip(n6823), .ck(clk), .q(
        \cache_data_A[4][49] ) );
  dp_1 \cache_data_A_reg[4][50]  ( .ip(n6822), .ck(clk), .q(
        \cache_data_A[4][50] ) );
  dp_1 \cache_data_A_reg[4][51]  ( .ip(n6821), .ck(clk), .q(
        \cache_data_A[4][51] ) );
  dp_1 \cache_data_A_reg[4][52]  ( .ip(n6820), .ck(clk), .q(
        \cache_data_A[4][52] ) );
  dp_1 \cache_data_A_reg[4][53]  ( .ip(n6819), .ck(clk), .q(
        \cache_data_A[4][53] ) );
  dp_1 \cache_data_A_reg[4][54]  ( .ip(n6818), .ck(clk), .q(
        \cache_data_A[4][54] ) );
  dp_1 \cache_data_A_reg[4][55]  ( .ip(n6817), .ck(clk), .q(
        \cache_data_A[4][55] ) );
  dp_1 \cache_data_A_reg[4][56]  ( .ip(n6816), .ck(clk), .q(
        \cache_data_A[4][56] ) );
  dp_1 \cache_data_A_reg[4][57]  ( .ip(n6815), .ck(clk), .q(
        \cache_data_A[4][57] ) );
  dp_1 \cache_data_A_reg[4][58]  ( .ip(n6814), .ck(clk), .q(
        \cache_data_A[4][58] ) );
  dp_1 \cache_data_A_reg[4][59]  ( .ip(n6813), .ck(clk), .q(
        \cache_data_A[4][59] ) );
  dp_1 \cache_data_A_reg[4][60]  ( .ip(n6812), .ck(clk), .q(
        \cache_data_A[4][60] ) );
  dp_1 \cache_data_A_reg[4][61]  ( .ip(n6811), .ck(clk), .q(
        \cache_data_A[4][61] ) );
  dp_1 \cache_data_A_reg[4][62]  ( .ip(n6810), .ck(clk), .q(
        \cache_data_A[4][62] ) );
  dp_1 \cache_data_A_reg[4][63]  ( .ip(n6809), .ck(clk), .q(
        \cache_data_A[4][63] ) );
  dp_1 \cache_data_A_reg[5][32]  ( .ip(n6712), .ck(clk), .q(
        \cache_data_A[5][32] ) );
  dp_1 \cache_data_A_reg[5][33]  ( .ip(n6711), .ck(clk), .q(
        \cache_data_A[5][33] ) );
  dp_1 \cache_data_A_reg[5][34]  ( .ip(n6710), .ck(clk), .q(
        \cache_data_A[5][34] ) );
  dp_1 \cache_data_A_reg[5][35]  ( .ip(n6709), .ck(clk), .q(
        \cache_data_A[5][35] ) );
  dp_1 \cache_data_A_reg[5][36]  ( .ip(n6708), .ck(clk), .q(
        \cache_data_A[5][36] ) );
  dp_1 \cache_data_A_reg[5][37]  ( .ip(n6707), .ck(clk), .q(
        \cache_data_A[5][37] ) );
  dp_1 \cache_data_A_reg[5][38]  ( .ip(n6706), .ck(clk), .q(
        \cache_data_A[5][38] ) );
  dp_1 \cache_data_A_reg[5][39]  ( .ip(n6705), .ck(clk), .q(
        \cache_data_A[5][39] ) );
  dp_1 \cache_data_A_reg[5][40]  ( .ip(n6704), .ck(clk), .q(
        \cache_data_A[5][40] ) );
  dp_1 \cache_data_A_reg[5][41]  ( .ip(n6703), .ck(clk), .q(
        \cache_data_A[5][41] ) );
  dp_1 \cache_data_A_reg[5][42]  ( .ip(n6702), .ck(clk), .q(
        \cache_data_A[5][42] ) );
  dp_1 \cache_data_A_reg[5][43]  ( .ip(n6701), .ck(clk), .q(
        \cache_data_A[5][43] ) );
  dp_1 \cache_data_A_reg[5][44]  ( .ip(n6700), .ck(clk), .q(
        \cache_data_A[5][44] ) );
  dp_1 \cache_data_A_reg[5][45]  ( .ip(n6699), .ck(clk), .q(
        \cache_data_A[5][45] ) );
  dp_1 \cache_data_A_reg[5][46]  ( .ip(n6698), .ck(clk), .q(
        \cache_data_A[5][46] ) );
  dp_1 \cache_data_A_reg[5][47]  ( .ip(n6697), .ck(clk), .q(
        \cache_data_A[5][47] ) );
  dp_1 \cache_data_A_reg[5][48]  ( .ip(n6696), .ck(clk), .q(
        \cache_data_A[5][48] ) );
  dp_1 \cache_data_A_reg[5][49]  ( .ip(n6695), .ck(clk), .q(
        \cache_data_A[5][49] ) );
  dp_1 \cache_data_A_reg[5][50]  ( .ip(n6694), .ck(clk), .q(
        \cache_data_A[5][50] ) );
  dp_1 \cache_data_A_reg[5][51]  ( .ip(n6693), .ck(clk), .q(
        \cache_data_A[5][51] ) );
  dp_1 \cache_data_A_reg[5][52]  ( .ip(n6692), .ck(clk), .q(
        \cache_data_A[5][52] ) );
  dp_1 \cache_data_A_reg[5][53]  ( .ip(n6691), .ck(clk), .q(
        \cache_data_A[5][53] ) );
  dp_1 \cache_data_A_reg[5][54]  ( .ip(n6690), .ck(clk), .q(
        \cache_data_A[5][54] ) );
  dp_1 \cache_data_A_reg[5][55]  ( .ip(n6689), .ck(clk), .q(
        \cache_data_A[5][55] ) );
  dp_1 \cache_data_A_reg[5][56]  ( .ip(n6688), .ck(clk), .q(
        \cache_data_A[5][56] ) );
  dp_1 \cache_data_A_reg[5][57]  ( .ip(n6687), .ck(clk), .q(
        \cache_data_A[5][57] ) );
  dp_1 \cache_data_A_reg[5][58]  ( .ip(n6686), .ck(clk), .q(
        \cache_data_A[5][58] ) );
  dp_1 \cache_data_A_reg[5][59]  ( .ip(n6685), .ck(clk), .q(
        \cache_data_A[5][59] ) );
  dp_1 \cache_data_A_reg[5][60]  ( .ip(n6684), .ck(clk), .q(
        \cache_data_A[5][60] ) );
  dp_1 \cache_data_A_reg[5][61]  ( .ip(n6683), .ck(clk), .q(
        \cache_data_A[5][61] ) );
  dp_1 \cache_data_A_reg[5][62]  ( .ip(n6682), .ck(clk), .q(
        \cache_data_A[5][62] ) );
  dp_1 \cache_data_A_reg[5][63]  ( .ip(n6681), .ck(clk), .q(
        \cache_data_A[5][63] ) );
  dp_1 \cache_data_A_reg[6][49]  ( .ip(n6584), .ck(clk), .q(
        \cache_data_A[6][49] ) );
  dp_1 \cache_data_A_reg[6][50]  ( .ip(n6583), .ck(clk), .q(
        \cache_data_A[6][50] ) );
  dp_1 \cache_data_A_reg[6][51]  ( .ip(n6582), .ck(clk), .q(
        \cache_data_A[6][51] ) );
  dp_1 \cache_data_A_reg[6][52]  ( .ip(n6581), .ck(clk), .q(
        \cache_data_A[6][52] ) );
  dp_1 \cache_data_A_reg[6][53]  ( .ip(n6580), .ck(clk), .q(
        \cache_data_A[6][53] ) );
  dp_1 \cache_data_A_reg[6][54]  ( .ip(n6579), .ck(clk), .q(
        \cache_data_A[6][54] ) );
  dp_1 \cache_data_A_reg[6][55]  ( .ip(n6578), .ck(clk), .q(
        \cache_data_A[6][55] ) );
  dp_1 \cache_data_A_reg[6][56]  ( .ip(n6577), .ck(clk), .q(
        \cache_data_A[6][56] ) );
  dp_1 \cache_data_A_reg[6][57]  ( .ip(n6576), .ck(clk), .q(
        \cache_data_A[6][57] ) );
  dp_1 \cache_data_A_reg[6][58]  ( .ip(n6575), .ck(clk), .q(
        \cache_data_A[6][58] ) );
  dp_1 \cache_data_A_reg[6][59]  ( .ip(n6574), .ck(clk), .q(
        \cache_data_A[6][59] ) );
  dp_1 \cache_data_A_reg[6][60]  ( .ip(n6573), .ck(clk), .q(
        \cache_data_A[6][60] ) );
  dp_1 \cache_data_A_reg[6][61]  ( .ip(n6572), .ck(clk), .q(
        \cache_data_A[6][61] ) );
  dp_1 \cache_data_A_reg[6][62]  ( .ip(n6571), .ck(clk), .q(
        \cache_data_A[6][62] ) );
  dp_1 \cache_data_A_reg[6][63]  ( .ip(n6570), .ck(clk), .q(
        \cache_data_A[6][63] ) );
  dp_1 \cache_data_A_reg[6][32]  ( .ip(n6569), .ck(clk), .q(
        \cache_data_A[6][32] ) );
  dp_1 \cache_data_A_reg[6][33]  ( .ip(n6568), .ck(clk), .q(
        \cache_data_A[6][33] ) );
  dp_1 \cache_data_A_reg[6][34]  ( .ip(n6567), .ck(clk), .q(
        \cache_data_A[6][34] ) );
  dp_1 \cache_data_A_reg[6][35]  ( .ip(n6566), .ck(clk), .q(
        \cache_data_A[6][35] ) );
  dp_1 \cache_data_A_reg[6][36]  ( .ip(n6565), .ck(clk), .q(
        \cache_data_A[6][36] ) );
  dp_1 \cache_data_A_reg[6][37]  ( .ip(n6564), .ck(clk), .q(
        \cache_data_A[6][37] ) );
  dp_1 \cache_data_A_reg[6][38]  ( .ip(n6563), .ck(clk), .q(
        \cache_data_A[6][38] ) );
  dp_1 \cache_data_A_reg[6][39]  ( .ip(n6562), .ck(clk), .q(
        \cache_data_A[6][39] ) );
  dp_1 \cache_data_A_reg[6][40]  ( .ip(n6561), .ck(clk), .q(
        \cache_data_A[6][40] ) );
  dp_1 \cache_data_A_reg[6][41]  ( .ip(n6560), .ck(clk), .q(
        \cache_data_A[6][41] ) );
  dp_1 \cache_data_A_reg[6][42]  ( .ip(n6559), .ck(clk), .q(
        \cache_data_A[6][42] ) );
  dp_1 \cache_data_A_reg[6][43]  ( .ip(n6558), .ck(clk), .q(
        \cache_data_A[6][43] ) );
  dp_1 \cache_data_A_reg[6][44]  ( .ip(n6557), .ck(clk), .q(
        \cache_data_A[6][44] ) );
  dp_1 \cache_data_A_reg[6][45]  ( .ip(n6556), .ck(clk), .q(
        \cache_data_A[6][45] ) );
  dp_1 \cache_data_A_reg[6][46]  ( .ip(n6555), .ck(clk), .q(
        \cache_data_A[6][46] ) );
  dp_1 \cache_data_A_reg[6][47]  ( .ip(n6554), .ck(clk), .q(
        \cache_data_A[6][47] ) );
  dp_1 \cache_data_A_reg[6][48]  ( .ip(n6553), .ck(clk), .q(
        \cache_data_A[6][48] ) );
  dp_1 \cache_data_A_reg[7][32]  ( .ip(n6456), .ck(clk), .q(
        \cache_data_A[7][32] ) );
  dp_1 \cache_data_A_reg[7][33]  ( .ip(n6455), .ck(clk), .q(
        \cache_data_A[7][33] ) );
  dp_1 \cache_data_A_reg[7][34]  ( .ip(n6454), .ck(clk), .q(
        \cache_data_A[7][34] ) );
  dp_1 \cache_data_A_reg[7][35]  ( .ip(n6453), .ck(clk), .q(
        \cache_data_A[7][35] ) );
  dp_1 \cache_data_A_reg[7][36]  ( .ip(n6452), .ck(clk), .q(
        \cache_data_A[7][36] ) );
  dp_1 \cache_data_A_reg[7][37]  ( .ip(n6451), .ck(clk), .q(
        \cache_data_A[7][37] ) );
  dp_1 \cache_data_A_reg[7][38]  ( .ip(n6450), .ck(clk), .q(
        \cache_data_A[7][38] ) );
  dp_1 \cache_data_A_reg[7][39]  ( .ip(n6449), .ck(clk), .q(
        \cache_data_A[7][39] ) );
  dp_1 \cache_data_A_reg[7][40]  ( .ip(n6448), .ck(clk), .q(
        \cache_data_A[7][40] ) );
  dp_1 \cache_data_A_reg[7][41]  ( .ip(n6447), .ck(clk), .q(
        \cache_data_A[7][41] ) );
  dp_1 \cache_data_A_reg[7][42]  ( .ip(n6446), .ck(clk), .q(
        \cache_data_A[7][42] ) );
  dp_1 \cache_data_A_reg[7][43]  ( .ip(n6445), .ck(clk), .q(
        \cache_data_A[7][43] ) );
  dp_1 \cache_data_A_reg[7][44]  ( .ip(n6444), .ck(clk), .q(
        \cache_data_A[7][44] ) );
  dp_1 \cache_data_A_reg[7][45]  ( .ip(n6443), .ck(clk), .q(
        \cache_data_A[7][45] ) );
  dp_1 \cache_data_A_reg[7][46]  ( .ip(n6442), .ck(clk), .q(
        \cache_data_A[7][46] ) );
  dp_1 \cache_data_A_reg[7][47]  ( .ip(n6441), .ck(clk), .q(
        \cache_data_A[7][47] ) );
  dp_1 \cache_data_A_reg[7][48]  ( .ip(n6440), .ck(clk), .q(
        \cache_data_A[7][48] ) );
  dp_1 \cache_data_A_reg[7][49]  ( .ip(n6439), .ck(clk), .q(
        \cache_data_A[7][49] ) );
  dp_1 \cache_data_A_reg[7][50]  ( .ip(n6438), .ck(clk), .q(
        \cache_data_A[7][50] ) );
  dp_1 \cache_data_A_reg[7][51]  ( .ip(n6437), .ck(clk), .q(
        \cache_data_A[7][51] ) );
  dp_1 \cache_data_A_reg[7][52]  ( .ip(n6436), .ck(clk), .q(
        \cache_data_A[7][52] ) );
  dp_1 \cache_data_A_reg[7][53]  ( .ip(n6435), .ck(clk), .q(
        \cache_data_A[7][53] ) );
  dp_1 \cache_data_A_reg[7][54]  ( .ip(n6434), .ck(clk), .q(
        \cache_data_A[7][54] ) );
  dp_1 \cache_data_A_reg[7][55]  ( .ip(n6433), .ck(clk), .q(
        \cache_data_A[7][55] ) );
  dp_1 \cache_data_A_reg[7][56]  ( .ip(n6432), .ck(clk), .q(
        \cache_data_A[7][56] ) );
  dp_1 \cache_data_A_reg[7][57]  ( .ip(n6431), .ck(clk), .q(
        \cache_data_A[7][57] ) );
  dp_1 \cache_data_A_reg[7][58]  ( .ip(n6430), .ck(clk), .q(
        \cache_data_A[7][58] ) );
  dp_1 \cache_data_A_reg[7][59]  ( .ip(n6429), .ck(clk), .q(
        \cache_data_A[7][59] ) );
  dp_1 \cache_data_A_reg[7][60]  ( .ip(n6428), .ck(clk), .q(
        \cache_data_A[7][60] ) );
  dp_1 \cache_data_A_reg[7][61]  ( .ip(n6427), .ck(clk), .q(
        \cache_data_A[7][61] ) );
  dp_1 \cache_data_A_reg[7][62]  ( .ip(n6426), .ck(clk), .q(
        \cache_data_A[7][62] ) );
  dp_1 \cache_data_A_reg[7][63]  ( .ip(n6425), .ck(clk), .q(
        \cache_data_A[7][63] ) );
  dp_1 \cache_data_A_reg[0][64]  ( .ip(n7320), .ck(clk), .q(
        \cache_data_A[0][64] ) );
  dp_1 \cache_data_A_reg[0][65]  ( .ip(n7319), .ck(clk), .q(
        \cache_data_A[0][65] ) );
  dp_1 \cache_data_A_reg[0][66]  ( .ip(n7318), .ck(clk), .q(
        \cache_data_A[0][66] ) );
  dp_1 \cache_data_A_reg[0][67]  ( .ip(n7317), .ck(clk), .q(
        \cache_data_A[0][67] ) );
  dp_1 \cache_data_A_reg[0][68]  ( .ip(n7316), .ck(clk), .q(
        \cache_data_A[0][68] ) );
  dp_1 \cache_data_A_reg[0][69]  ( .ip(n7315), .ck(clk), .q(
        \cache_data_A[0][69] ) );
  dp_1 \cache_data_A_reg[0][70]  ( .ip(n7314), .ck(clk), .q(
        \cache_data_A[0][70] ) );
  dp_1 \cache_data_A_reg[0][71]  ( .ip(n7313), .ck(clk), .q(
        \cache_data_A[0][71] ) );
  dp_1 \cache_data_A_reg[0][72]  ( .ip(n7312), .ck(clk), .q(
        \cache_data_A[0][72] ) );
  dp_1 \cache_data_A_reg[0][73]  ( .ip(n7311), .ck(clk), .q(
        \cache_data_A[0][73] ) );
  dp_1 \cache_data_A_reg[0][74]  ( .ip(n7310), .ck(clk), .q(
        \cache_data_A[0][74] ) );
  dp_1 \cache_data_A_reg[0][75]  ( .ip(n7309), .ck(clk), .q(
        \cache_data_A[0][75] ) );
  dp_1 \cache_data_A_reg[0][76]  ( .ip(n7308), .ck(clk), .q(
        \cache_data_A[0][76] ) );
  dp_1 \cache_data_A_reg[0][77]  ( .ip(n7307), .ck(clk), .q(
        \cache_data_A[0][77] ) );
  dp_1 \cache_data_A_reg[0][78]  ( .ip(n7306), .ck(clk), .q(
        \cache_data_A[0][78] ) );
  dp_1 \cache_data_A_reg[0][79]  ( .ip(n7305), .ck(clk), .q(
        \cache_data_A[0][79] ) );
  dp_1 \cache_data_A_reg[0][80]  ( .ip(n7304), .ck(clk), .q(
        \cache_data_A[0][80] ) );
  dp_1 \cache_data_A_reg[0][81]  ( .ip(n7303), .ck(clk), .q(
        \cache_data_A[0][81] ) );
  dp_1 \cache_data_A_reg[0][82]  ( .ip(n7302), .ck(clk), .q(
        \cache_data_A[0][82] ) );
  dp_1 \cache_data_A_reg[0][83]  ( .ip(n7301), .ck(clk), .q(
        \cache_data_A[0][83] ) );
  dp_1 \cache_data_A_reg[0][84]  ( .ip(n7300), .ck(clk), .q(
        \cache_data_A[0][84] ) );
  dp_1 \cache_data_A_reg[0][85]  ( .ip(n7299), .ck(clk), .q(
        \cache_data_A[0][85] ) );
  dp_1 \cache_data_A_reg[0][86]  ( .ip(n7298), .ck(clk), .q(
        \cache_data_A[0][86] ) );
  dp_1 \cache_data_A_reg[0][87]  ( .ip(n7297), .ck(clk), .q(
        \cache_data_A[0][87] ) );
  dp_1 \cache_data_A_reg[0][88]  ( .ip(n7296), .ck(clk), .q(
        \cache_data_A[0][88] ) );
  dp_1 \cache_data_A_reg[0][89]  ( .ip(n7295), .ck(clk), .q(
        \cache_data_A[0][89] ) );
  dp_1 \cache_data_A_reg[0][90]  ( .ip(n7294), .ck(clk), .q(
        \cache_data_A[0][90] ) );
  dp_1 \cache_data_A_reg[0][91]  ( .ip(n7293), .ck(clk), .q(
        \cache_data_A[0][91] ) );
  dp_1 \cache_data_A_reg[0][92]  ( .ip(n7292), .ck(clk), .q(
        \cache_data_A[0][92] ) );
  dp_1 \cache_data_A_reg[0][93]  ( .ip(n7291), .ck(clk), .q(
        \cache_data_A[0][93] ) );
  dp_1 \cache_data_A_reg[0][94]  ( .ip(n7290), .ck(clk), .q(
        \cache_data_A[0][94] ) );
  dp_1 \cache_data_A_reg[0][95]  ( .ip(n7289), .ck(clk), .q(
        \cache_data_A[0][95] ) );
  dp_1 \cache_data_A_reg[1][95]  ( .ip(n7192), .ck(clk), .q(
        \cache_data_A[1][95] ) );
  dp_1 \cache_data_A_reg[1][64]  ( .ip(n7191), .ck(clk), .q(
        \cache_data_A[1][64] ) );
  dp_1 \cache_data_A_reg[1][65]  ( .ip(n7190), .ck(clk), .q(
        \cache_data_A[1][65] ) );
  dp_1 \cache_data_A_reg[1][66]  ( .ip(n7189), .ck(clk), .q(
        \cache_data_A[1][66] ) );
  dp_1 \cache_data_A_reg[1][67]  ( .ip(n7188), .ck(clk), .q(
        \cache_data_A[1][67] ) );
  dp_1 \cache_data_A_reg[1][68]  ( .ip(n7187), .ck(clk), .q(
        \cache_data_A[1][68] ) );
  dp_1 \cache_data_A_reg[1][69]  ( .ip(n7186), .ck(clk), .q(
        \cache_data_A[1][69] ) );
  dp_1 \cache_data_A_reg[1][70]  ( .ip(n7185), .ck(clk), .q(
        \cache_data_A[1][70] ) );
  dp_1 \cache_data_A_reg[1][71]  ( .ip(n7184), .ck(clk), .q(
        \cache_data_A[1][71] ) );
  dp_1 \cache_data_A_reg[1][72]  ( .ip(n7183), .ck(clk), .q(
        \cache_data_A[1][72] ) );
  dp_1 \cache_data_A_reg[1][73]  ( .ip(n7182), .ck(clk), .q(
        \cache_data_A[1][73] ) );
  dp_1 \cache_data_A_reg[1][74]  ( .ip(n7181), .ck(clk), .q(
        \cache_data_A[1][74] ) );
  dp_1 \cache_data_A_reg[1][75]  ( .ip(n7180), .ck(clk), .q(
        \cache_data_A[1][75] ) );
  dp_1 \cache_data_A_reg[1][76]  ( .ip(n7179), .ck(clk), .q(
        \cache_data_A[1][76] ) );
  dp_1 \cache_data_A_reg[1][77]  ( .ip(n7178), .ck(clk), .q(
        \cache_data_A[1][77] ) );
  dp_1 \cache_data_A_reg[1][78]  ( .ip(n7177), .ck(clk), .q(
        \cache_data_A[1][78] ) );
  dp_1 \cache_data_A_reg[1][79]  ( .ip(n7176), .ck(clk), .q(
        \cache_data_A[1][79] ) );
  dp_1 \cache_data_A_reg[1][80]  ( .ip(n7175), .ck(clk), .q(
        \cache_data_A[1][80] ) );
  dp_1 \cache_data_A_reg[1][81]  ( .ip(n7174), .ck(clk), .q(
        \cache_data_A[1][81] ) );
  dp_1 \cache_data_A_reg[1][82]  ( .ip(n7173), .ck(clk), .q(
        \cache_data_A[1][82] ) );
  dp_1 \cache_data_A_reg[1][83]  ( .ip(n7172), .ck(clk), .q(
        \cache_data_A[1][83] ) );
  dp_1 \cache_data_A_reg[1][84]  ( .ip(n7171), .ck(clk), .q(
        \cache_data_A[1][84] ) );
  dp_1 \cache_data_A_reg[1][85]  ( .ip(n7170), .ck(clk), .q(
        \cache_data_A[1][85] ) );
  dp_1 \cache_data_A_reg[1][86]  ( .ip(n7169), .ck(clk), .q(
        \cache_data_A[1][86] ) );
  dp_1 \cache_data_A_reg[1][87]  ( .ip(n7168), .ck(clk), .q(
        \cache_data_A[1][87] ) );
  dp_1 \cache_data_A_reg[1][88]  ( .ip(n7167), .ck(clk), .q(
        \cache_data_A[1][88] ) );
  dp_1 \cache_data_A_reg[1][89]  ( .ip(n7166), .ck(clk), .q(
        \cache_data_A[1][89] ) );
  dp_1 \cache_data_A_reg[1][90]  ( .ip(n7165), .ck(clk), .q(
        \cache_data_A[1][90] ) );
  dp_1 \cache_data_A_reg[1][91]  ( .ip(n7164), .ck(clk), .q(
        \cache_data_A[1][91] ) );
  dp_1 \cache_data_A_reg[1][92]  ( .ip(n7163), .ck(clk), .q(
        \cache_data_A[1][92] ) );
  dp_1 \cache_data_A_reg[1][93]  ( .ip(n7162), .ck(clk), .q(
        \cache_data_A[1][93] ) );
  dp_1 \cache_data_A_reg[1][94]  ( .ip(n7161), .ck(clk), .q(
        \cache_data_A[1][94] ) );
  dp_1 \cache_data_A_reg[2][66]  ( .ip(n7064), .ck(clk), .q(
        \cache_data_A[2][66] ) );
  dp_1 \cache_data_A_reg[2][67]  ( .ip(n7063), .ck(clk), .q(
        \cache_data_A[2][67] ) );
  dp_1 \cache_data_A_reg[2][68]  ( .ip(n7062), .ck(clk), .q(
        \cache_data_A[2][68] ) );
  dp_1 \cache_data_A_reg[2][69]  ( .ip(n7061), .ck(clk), .q(
        \cache_data_A[2][69] ) );
  dp_1 \cache_data_A_reg[2][70]  ( .ip(n7060), .ck(clk), .q(
        \cache_data_A[2][70] ) );
  dp_1 \cache_data_A_reg[2][71]  ( .ip(n7059), .ck(clk), .q(
        \cache_data_A[2][71] ) );
  dp_1 \cache_data_A_reg[2][72]  ( .ip(n7058), .ck(clk), .q(
        \cache_data_A[2][72] ) );
  dp_1 \cache_data_A_reg[2][73]  ( .ip(n7057), .ck(clk), .q(
        \cache_data_A[2][73] ) );
  dp_1 \cache_data_A_reg[2][74]  ( .ip(n7056), .ck(clk), .q(
        \cache_data_A[2][74] ) );
  dp_1 \cache_data_A_reg[2][75]  ( .ip(n7055), .ck(clk), .q(
        \cache_data_A[2][75] ) );
  dp_1 \cache_data_A_reg[2][76]  ( .ip(n7054), .ck(clk), .q(
        \cache_data_A[2][76] ) );
  dp_1 \cache_data_A_reg[2][77]  ( .ip(n7053), .ck(clk), .q(
        \cache_data_A[2][77] ) );
  dp_1 \cache_data_A_reg[2][78]  ( .ip(n7052), .ck(clk), .q(
        \cache_data_A[2][78] ) );
  dp_1 \cache_data_A_reg[2][79]  ( .ip(n7051), .ck(clk), .q(
        \cache_data_A[2][79] ) );
  dp_1 \cache_data_A_reg[2][80]  ( .ip(n7050), .ck(clk), .q(
        \cache_data_A[2][80] ) );
  dp_1 \cache_data_A_reg[2][81]  ( .ip(n7049), .ck(clk), .q(
        \cache_data_A[2][81] ) );
  dp_1 \cache_data_A_reg[2][82]  ( .ip(n7048), .ck(clk), .q(
        \cache_data_A[2][82] ) );
  dp_1 \cache_data_A_reg[2][83]  ( .ip(n7047), .ck(clk), .q(
        \cache_data_A[2][83] ) );
  dp_1 \cache_data_A_reg[2][84]  ( .ip(n7046), .ck(clk), .q(
        \cache_data_A[2][84] ) );
  dp_1 \cache_data_A_reg[2][85]  ( .ip(n7045), .ck(clk), .q(
        \cache_data_A[2][85] ) );
  dp_1 \cache_data_A_reg[2][86]  ( .ip(n7044), .ck(clk), .q(
        \cache_data_A[2][86] ) );
  dp_1 \cache_data_A_reg[2][87]  ( .ip(n7043), .ck(clk), .q(
        \cache_data_A[2][87] ) );
  dp_1 \cache_data_A_reg[2][88]  ( .ip(n7042), .ck(clk), .q(
        \cache_data_A[2][88] ) );
  dp_1 \cache_data_A_reg[2][89]  ( .ip(n7041), .ck(clk), .q(
        \cache_data_A[2][89] ) );
  dp_1 \cache_data_A_reg[2][90]  ( .ip(n7040), .ck(clk), .q(
        \cache_data_A[2][90] ) );
  dp_1 \cache_data_A_reg[2][91]  ( .ip(n7039), .ck(clk), .q(
        \cache_data_A[2][91] ) );
  dp_1 \cache_data_A_reg[2][92]  ( .ip(n7038), .ck(clk), .q(
        \cache_data_A[2][92] ) );
  dp_1 \cache_data_A_reg[2][93]  ( .ip(n7037), .ck(clk), .q(
        \cache_data_A[2][93] ) );
  dp_1 \cache_data_A_reg[2][94]  ( .ip(n7036), .ck(clk), .q(
        \cache_data_A[2][94] ) );
  dp_1 \cache_data_A_reg[2][95]  ( .ip(n7035), .ck(clk), .q(
        \cache_data_A[2][95] ) );
  dp_1 \cache_data_A_reg[2][64]  ( .ip(n7034), .ck(clk), .q(
        \cache_data_A[2][64] ) );
  dp_1 \cache_data_A_reg[2][65]  ( .ip(n7033), .ck(clk), .q(
        \cache_data_A[2][65] ) );
  dp_1 \cache_data_A_reg[3][64]  ( .ip(n6936), .ck(clk), .q(
        \cache_data_A[3][64] ) );
  dp_1 \cache_data_A_reg[3][65]  ( .ip(n6935), .ck(clk), .q(
        \cache_data_A[3][65] ) );
  dp_1 \cache_data_A_reg[3][66]  ( .ip(n6934), .ck(clk), .q(
        \cache_data_A[3][66] ) );
  dp_1 \cache_data_A_reg[3][67]  ( .ip(n6933), .ck(clk), .q(
        \cache_data_A[3][67] ) );
  dp_1 \cache_data_A_reg[3][68]  ( .ip(n6932), .ck(clk), .q(
        \cache_data_A[3][68] ) );
  dp_1 \cache_data_A_reg[3][69]  ( .ip(n6931), .ck(clk), .q(
        \cache_data_A[3][69] ) );
  dp_1 \cache_data_A_reg[3][70]  ( .ip(n6930), .ck(clk), .q(
        \cache_data_A[3][70] ) );
  dp_1 \cache_data_A_reg[3][71]  ( .ip(n6929), .ck(clk), .q(
        \cache_data_A[3][71] ) );
  dp_1 \cache_data_A_reg[3][72]  ( .ip(n6928), .ck(clk), .q(
        \cache_data_A[3][72] ) );
  dp_1 \cache_data_A_reg[3][73]  ( .ip(n6927), .ck(clk), .q(
        \cache_data_A[3][73] ) );
  dp_1 \cache_data_A_reg[3][74]  ( .ip(n6926), .ck(clk), .q(
        \cache_data_A[3][74] ) );
  dp_1 \cache_data_A_reg[3][75]  ( .ip(n6925), .ck(clk), .q(
        \cache_data_A[3][75] ) );
  dp_1 \cache_data_A_reg[3][76]  ( .ip(n6924), .ck(clk), .q(
        \cache_data_A[3][76] ) );
  dp_1 \cache_data_A_reg[3][77]  ( .ip(n6923), .ck(clk), .q(
        \cache_data_A[3][77] ) );
  dp_1 \cache_data_A_reg[3][78]  ( .ip(n6922), .ck(clk), .q(
        \cache_data_A[3][78] ) );
  dp_1 \cache_data_A_reg[3][79]  ( .ip(n6921), .ck(clk), .q(
        \cache_data_A[3][79] ) );
  dp_1 \cache_data_A_reg[3][80]  ( .ip(n6920), .ck(clk), .q(
        \cache_data_A[3][80] ) );
  dp_1 \cache_data_A_reg[3][81]  ( .ip(n6919), .ck(clk), .q(
        \cache_data_A[3][81] ) );
  dp_1 \cache_data_A_reg[3][82]  ( .ip(n6918), .ck(clk), .q(
        \cache_data_A[3][82] ) );
  dp_1 \cache_data_A_reg[3][83]  ( .ip(n6917), .ck(clk), .q(
        \cache_data_A[3][83] ) );
  dp_1 \cache_data_A_reg[3][84]  ( .ip(n6916), .ck(clk), .q(
        \cache_data_A[3][84] ) );
  dp_1 \cache_data_A_reg[3][85]  ( .ip(n6915), .ck(clk), .q(
        \cache_data_A[3][85] ) );
  dp_1 \cache_data_A_reg[3][86]  ( .ip(n6914), .ck(clk), .q(
        \cache_data_A[3][86] ) );
  dp_1 \cache_data_A_reg[3][87]  ( .ip(n6913), .ck(clk), .q(
        \cache_data_A[3][87] ) );
  dp_1 \cache_data_A_reg[3][88]  ( .ip(n6912), .ck(clk), .q(
        \cache_data_A[3][88] ) );
  dp_1 \cache_data_A_reg[3][89]  ( .ip(n6911), .ck(clk), .q(
        \cache_data_A[3][89] ) );
  dp_1 \cache_data_A_reg[3][90]  ( .ip(n6910), .ck(clk), .q(
        \cache_data_A[3][90] ) );
  dp_1 \cache_data_A_reg[3][91]  ( .ip(n6909), .ck(clk), .q(
        \cache_data_A[3][91] ) );
  dp_1 \cache_data_A_reg[3][92]  ( .ip(n6908), .ck(clk), .q(
        \cache_data_A[3][92] ) );
  dp_1 \cache_data_A_reg[3][93]  ( .ip(n6907), .ck(clk), .q(
        \cache_data_A[3][93] ) );
  dp_1 \cache_data_A_reg[3][94]  ( .ip(n6906), .ck(clk), .q(
        \cache_data_A[3][94] ) );
  dp_1 \cache_data_A_reg[3][95]  ( .ip(n6905), .ck(clk), .q(
        \cache_data_A[3][95] ) );
  dp_1 \cache_data_A_reg[4][64]  ( .ip(n6808), .ck(clk), .q(
        \cache_data_A[4][64] ) );
  dp_1 \cache_data_A_reg[4][65]  ( .ip(n6807), .ck(clk), .q(
        \cache_data_A[4][65] ) );
  dp_1 \cache_data_A_reg[4][66]  ( .ip(n6806), .ck(clk), .q(
        \cache_data_A[4][66] ) );
  dp_1 \cache_data_A_reg[4][67]  ( .ip(n6805), .ck(clk), .q(
        \cache_data_A[4][67] ) );
  dp_1 \cache_data_A_reg[4][68]  ( .ip(n6804), .ck(clk), .q(
        \cache_data_A[4][68] ) );
  dp_1 \cache_data_A_reg[4][69]  ( .ip(n6803), .ck(clk), .q(
        \cache_data_A[4][69] ) );
  dp_1 \cache_data_A_reg[4][70]  ( .ip(n6802), .ck(clk), .q(
        \cache_data_A[4][70] ) );
  dp_1 \cache_data_A_reg[4][71]  ( .ip(n6801), .ck(clk), .q(
        \cache_data_A[4][71] ) );
  dp_1 \cache_data_A_reg[4][72]  ( .ip(n6800), .ck(clk), .q(
        \cache_data_A[4][72] ) );
  dp_1 \cache_data_A_reg[4][73]  ( .ip(n6799), .ck(clk), .q(
        \cache_data_A[4][73] ) );
  dp_1 \cache_data_A_reg[4][74]  ( .ip(n6798), .ck(clk), .q(
        \cache_data_A[4][74] ) );
  dp_1 \cache_data_A_reg[4][75]  ( .ip(n6797), .ck(clk), .q(
        \cache_data_A[4][75] ) );
  dp_1 \cache_data_A_reg[4][76]  ( .ip(n6796), .ck(clk), .q(
        \cache_data_A[4][76] ) );
  dp_1 \cache_data_A_reg[4][77]  ( .ip(n6795), .ck(clk), .q(
        \cache_data_A[4][77] ) );
  dp_1 \cache_data_A_reg[4][78]  ( .ip(n6794), .ck(clk), .q(
        \cache_data_A[4][78] ) );
  dp_1 \cache_data_A_reg[4][79]  ( .ip(n6793), .ck(clk), .q(
        \cache_data_A[4][79] ) );
  dp_1 \cache_data_A_reg[4][80]  ( .ip(n6792), .ck(clk), .q(
        \cache_data_A[4][80] ) );
  dp_1 \cache_data_A_reg[4][81]  ( .ip(n6791), .ck(clk), .q(
        \cache_data_A[4][81] ) );
  dp_1 \cache_data_A_reg[4][82]  ( .ip(n6790), .ck(clk), .q(
        \cache_data_A[4][82] ) );
  dp_1 \cache_data_A_reg[4][83]  ( .ip(n6789), .ck(clk), .q(
        \cache_data_A[4][83] ) );
  dp_1 \cache_data_A_reg[4][84]  ( .ip(n6788), .ck(clk), .q(
        \cache_data_A[4][84] ) );
  dp_1 \cache_data_A_reg[4][85]  ( .ip(n6787), .ck(clk), .q(
        \cache_data_A[4][85] ) );
  dp_1 \cache_data_A_reg[4][86]  ( .ip(n6786), .ck(clk), .q(
        \cache_data_A[4][86] ) );
  dp_1 \cache_data_A_reg[4][87]  ( .ip(n6785), .ck(clk), .q(
        \cache_data_A[4][87] ) );
  dp_1 \cache_data_A_reg[4][88]  ( .ip(n6784), .ck(clk), .q(
        \cache_data_A[4][88] ) );
  dp_1 \cache_data_A_reg[4][89]  ( .ip(n6783), .ck(clk), .q(
        \cache_data_A[4][89] ) );
  dp_1 \cache_data_A_reg[4][90]  ( .ip(n6782), .ck(clk), .q(
        \cache_data_A[4][90] ) );
  dp_1 \cache_data_A_reg[4][91]  ( .ip(n6781), .ck(clk), .q(
        \cache_data_A[4][91] ) );
  dp_1 \cache_data_A_reg[4][92]  ( .ip(n6780), .ck(clk), .q(
        \cache_data_A[4][92] ) );
  dp_1 \cache_data_A_reg[4][93]  ( .ip(n6779), .ck(clk), .q(
        \cache_data_A[4][93] ) );
  dp_1 \cache_data_A_reg[4][94]  ( .ip(n6778), .ck(clk), .q(
        \cache_data_A[4][94] ) );
  dp_1 \cache_data_A_reg[4][95]  ( .ip(n6777), .ck(clk), .q(
        \cache_data_A[4][95] ) );
  dp_1 \cache_data_A_reg[5][78]  ( .ip(n6680), .ck(clk), .q(
        \cache_data_A[5][78] ) );
  dp_1 \cache_data_A_reg[5][79]  ( .ip(n6679), .ck(clk), .q(
        \cache_data_A[5][79] ) );
  dp_1 \cache_data_A_reg[5][80]  ( .ip(n6678), .ck(clk), .q(
        \cache_data_A[5][80] ) );
  dp_1 \cache_data_A_reg[5][81]  ( .ip(n6677), .ck(clk), .q(
        \cache_data_A[5][81] ) );
  dp_1 \cache_data_A_reg[5][82]  ( .ip(n6676), .ck(clk), .q(
        \cache_data_A[5][82] ) );
  dp_1 \cache_data_A_reg[5][83]  ( .ip(n6675), .ck(clk), .q(
        \cache_data_A[5][83] ) );
  dp_1 \cache_data_A_reg[5][84]  ( .ip(n6674), .ck(clk), .q(
        \cache_data_A[5][84] ) );
  dp_1 \cache_data_A_reg[5][85]  ( .ip(n6673), .ck(clk), .q(
        \cache_data_A[5][85] ) );
  dp_1 \cache_data_A_reg[5][86]  ( .ip(n6672), .ck(clk), .q(
        \cache_data_A[5][86] ) );
  dp_1 \cache_data_A_reg[5][87]  ( .ip(n6671), .ck(clk), .q(
        \cache_data_A[5][87] ) );
  dp_1 \cache_data_A_reg[5][88]  ( .ip(n6670), .ck(clk), .q(
        \cache_data_A[5][88] ) );
  dp_1 \cache_data_A_reg[5][89]  ( .ip(n6669), .ck(clk), .q(
        \cache_data_A[5][89] ) );
  dp_1 \cache_data_A_reg[5][90]  ( .ip(n6668), .ck(clk), .q(
        \cache_data_A[5][90] ) );
  dp_1 \cache_data_A_reg[5][91]  ( .ip(n6667), .ck(clk), .q(
        \cache_data_A[5][91] ) );
  dp_1 \cache_data_A_reg[5][92]  ( .ip(n6666), .ck(clk), .q(
        \cache_data_A[5][92] ) );
  dp_1 \cache_data_A_reg[5][93]  ( .ip(n6665), .ck(clk), .q(
        \cache_data_A[5][93] ) );
  dp_1 \cache_data_A_reg[5][94]  ( .ip(n6664), .ck(clk), .q(
        \cache_data_A[5][94] ) );
  dp_1 \cache_data_A_reg[5][95]  ( .ip(n6663), .ck(clk), .q(
        \cache_data_A[5][95] ) );
  dp_1 \cache_data_A_reg[5][64]  ( .ip(n6662), .ck(clk), .q(
        \cache_data_A[5][64] ) );
  dp_1 \cache_data_A_reg[5][65]  ( .ip(n6661), .ck(clk), .q(
        \cache_data_A[5][65] ) );
  dp_1 \cache_data_A_reg[5][66]  ( .ip(n6660), .ck(clk), .q(
        \cache_data_A[5][66] ) );
  dp_1 \cache_data_A_reg[5][67]  ( .ip(n6659), .ck(clk), .q(
        \cache_data_A[5][67] ) );
  dp_1 \cache_data_A_reg[5][68]  ( .ip(n6658), .ck(clk), .q(
        \cache_data_A[5][68] ) );
  dp_1 \cache_data_A_reg[5][69]  ( .ip(n6657), .ck(clk), .q(
        \cache_data_A[5][69] ) );
  dp_1 \cache_data_A_reg[5][70]  ( .ip(n6656), .ck(clk), .q(
        \cache_data_A[5][70] ) );
  dp_1 \cache_data_A_reg[5][71]  ( .ip(n6655), .ck(clk), .q(
        \cache_data_A[5][71] ) );
  dp_1 \cache_data_A_reg[5][72]  ( .ip(n6654), .ck(clk), .q(
        \cache_data_A[5][72] ) );
  dp_1 \cache_data_A_reg[5][73]  ( .ip(n6653), .ck(clk), .q(
        \cache_data_A[5][73] ) );
  dp_1 \cache_data_A_reg[5][74]  ( .ip(n6652), .ck(clk), .q(
        \cache_data_A[5][74] ) );
  dp_1 \cache_data_A_reg[5][75]  ( .ip(n6651), .ck(clk), .q(
        \cache_data_A[5][75] ) );
  dp_1 \cache_data_A_reg[5][76]  ( .ip(n6650), .ck(clk), .q(
        \cache_data_A[5][76] ) );
  dp_1 \cache_data_A_reg[5][77]  ( .ip(n6649), .ck(clk), .q(
        \cache_data_A[5][77] ) );
  dp_1 \cache_data_A_reg[6][64]  ( .ip(n6552), .ck(clk), .q(
        \cache_data_A[6][64] ) );
  dp_1 \cache_data_A_reg[6][65]  ( .ip(n6551), .ck(clk), .q(
        \cache_data_A[6][65] ) );
  dp_1 \cache_data_A_reg[6][66]  ( .ip(n6550), .ck(clk), .q(
        \cache_data_A[6][66] ) );
  dp_1 \cache_data_A_reg[6][67]  ( .ip(n6549), .ck(clk), .q(
        \cache_data_A[6][67] ) );
  dp_1 \cache_data_A_reg[6][68]  ( .ip(n6548), .ck(clk), .q(
        \cache_data_A[6][68] ) );
  dp_1 \cache_data_A_reg[6][69]  ( .ip(n6547), .ck(clk), .q(
        \cache_data_A[6][69] ) );
  dp_1 \cache_data_A_reg[6][70]  ( .ip(n6546), .ck(clk), .q(
        \cache_data_A[6][70] ) );
  dp_1 \cache_data_A_reg[6][71]  ( .ip(n6545), .ck(clk), .q(
        \cache_data_A[6][71] ) );
  dp_1 \cache_data_A_reg[6][72]  ( .ip(n6544), .ck(clk), .q(
        \cache_data_A[6][72] ) );
  dp_1 \cache_data_A_reg[6][73]  ( .ip(n6543), .ck(clk), .q(
        \cache_data_A[6][73] ) );
  dp_1 \cache_data_A_reg[6][74]  ( .ip(n6542), .ck(clk), .q(
        \cache_data_A[6][74] ) );
  dp_1 \cache_data_A_reg[6][75]  ( .ip(n6541), .ck(clk), .q(
        \cache_data_A[6][75] ) );
  dp_1 \cache_data_A_reg[6][76]  ( .ip(n6540), .ck(clk), .q(
        \cache_data_A[6][76] ) );
  dp_1 \cache_data_A_reg[6][77]  ( .ip(n6539), .ck(clk), .q(
        \cache_data_A[6][77] ) );
  dp_1 \cache_data_A_reg[6][78]  ( .ip(n6538), .ck(clk), .q(
        \cache_data_A[6][78] ) );
  dp_1 \cache_data_A_reg[6][79]  ( .ip(n6537), .ck(clk), .q(
        \cache_data_A[6][79] ) );
  dp_1 \cache_data_A_reg[6][80]  ( .ip(n6536), .ck(clk), .q(
        \cache_data_A[6][80] ) );
  dp_1 \cache_data_A_reg[6][81]  ( .ip(n6535), .ck(clk), .q(
        \cache_data_A[6][81] ) );
  dp_1 \cache_data_A_reg[6][82]  ( .ip(n6534), .ck(clk), .q(
        \cache_data_A[6][82] ) );
  dp_1 \cache_data_A_reg[6][83]  ( .ip(n6533), .ck(clk), .q(
        \cache_data_A[6][83] ) );
  dp_1 \cache_data_A_reg[6][84]  ( .ip(n6532), .ck(clk), .q(
        \cache_data_A[6][84] ) );
  dp_1 \cache_data_A_reg[6][85]  ( .ip(n6531), .ck(clk), .q(
        \cache_data_A[6][85] ) );
  dp_1 \cache_data_A_reg[6][86]  ( .ip(n6530), .ck(clk), .q(
        \cache_data_A[6][86] ) );
  dp_1 \cache_data_A_reg[6][87]  ( .ip(n6529), .ck(clk), .q(
        \cache_data_A[6][87] ) );
  dp_1 \cache_data_A_reg[6][88]  ( .ip(n6528), .ck(clk), .q(
        \cache_data_A[6][88] ) );
  dp_1 \cache_data_A_reg[6][89]  ( .ip(n6527), .ck(clk), .q(
        \cache_data_A[6][89] ) );
  dp_1 \cache_data_A_reg[6][90]  ( .ip(n6526), .ck(clk), .q(
        \cache_data_A[6][90] ) );
  dp_1 \cache_data_A_reg[6][91]  ( .ip(n6525), .ck(clk), .q(
        \cache_data_A[6][91] ) );
  dp_1 \cache_data_A_reg[6][92]  ( .ip(n6524), .ck(clk), .q(
        \cache_data_A[6][92] ) );
  dp_1 \cache_data_A_reg[6][93]  ( .ip(n6523), .ck(clk), .q(
        \cache_data_A[6][93] ) );
  dp_1 \cache_data_A_reg[6][94]  ( .ip(n6522), .ck(clk), .q(
        \cache_data_A[6][94] ) );
  dp_1 \cache_data_A_reg[6][95]  ( .ip(n6521), .ck(clk), .q(
        \cache_data_A[6][95] ) );
  dp_1 \cache_data_A_reg[7][64]  ( .ip(n6424), .ck(clk), .q(
        \cache_data_A[7][64] ) );
  dp_1 \cache_data_A_reg[7][65]  ( .ip(n6423), .ck(clk), .q(
        \cache_data_A[7][65] ) );
  dp_1 \cache_data_A_reg[7][66]  ( .ip(n6422), .ck(clk), .q(
        \cache_data_A[7][66] ) );
  dp_1 \cache_data_A_reg[7][67]  ( .ip(n6421), .ck(clk), .q(
        \cache_data_A[7][67] ) );
  dp_1 \cache_data_A_reg[7][68]  ( .ip(n6420), .ck(clk), .q(
        \cache_data_A[7][68] ) );
  dp_1 \cache_data_A_reg[7][69]  ( .ip(n6419), .ck(clk), .q(
        \cache_data_A[7][69] ) );
  dp_1 \cache_data_A_reg[7][70]  ( .ip(n6418), .ck(clk), .q(
        \cache_data_A[7][70] ) );
  dp_1 \cache_data_A_reg[7][71]  ( .ip(n6417), .ck(clk), .q(
        \cache_data_A[7][71] ) );
  dp_1 \cache_data_A_reg[7][72]  ( .ip(n6416), .ck(clk), .q(
        \cache_data_A[7][72] ) );
  dp_1 \cache_data_A_reg[7][73]  ( .ip(n6415), .ck(clk), .q(
        \cache_data_A[7][73] ) );
  dp_1 \cache_data_A_reg[7][74]  ( .ip(n6414), .ck(clk), .q(
        \cache_data_A[7][74] ) );
  dp_1 \cache_data_A_reg[7][75]  ( .ip(n6413), .ck(clk), .q(
        \cache_data_A[7][75] ) );
  dp_1 \cache_data_A_reg[7][76]  ( .ip(n6412), .ck(clk), .q(
        \cache_data_A[7][76] ) );
  dp_1 \cache_data_A_reg[7][77]  ( .ip(n6411), .ck(clk), .q(
        \cache_data_A[7][77] ) );
  dp_1 \cache_data_A_reg[7][78]  ( .ip(n6410), .ck(clk), .q(
        \cache_data_A[7][78] ) );
  dp_1 \cache_data_A_reg[7][79]  ( .ip(n6409), .ck(clk), .q(
        \cache_data_A[7][79] ) );
  dp_1 \cache_data_A_reg[7][80]  ( .ip(n6408), .ck(clk), .q(
        \cache_data_A[7][80] ) );
  dp_1 \cache_data_A_reg[7][81]  ( .ip(n6407), .ck(clk), .q(
        \cache_data_A[7][81] ) );
  dp_1 \cache_data_A_reg[7][82]  ( .ip(n6406), .ck(clk), .q(
        \cache_data_A[7][82] ) );
  dp_1 \cache_data_A_reg[7][83]  ( .ip(n6405), .ck(clk), .q(
        \cache_data_A[7][83] ) );
  dp_1 \cache_data_A_reg[7][84]  ( .ip(n6404), .ck(clk), .q(
        \cache_data_A[7][84] ) );
  dp_1 \cache_data_A_reg[7][85]  ( .ip(n6403), .ck(clk), .q(
        \cache_data_A[7][85] ) );
  dp_1 \cache_data_A_reg[7][86]  ( .ip(n6402), .ck(clk), .q(
        \cache_data_A[7][86] ) );
  dp_1 \cache_data_A_reg[7][87]  ( .ip(n6401), .ck(clk), .q(
        \cache_data_A[7][87] ) );
  dp_1 \cache_data_A_reg[7][88]  ( .ip(n6400), .ck(clk), .q(
        \cache_data_A[7][88] ) );
  dp_1 \cache_data_A_reg[7][89]  ( .ip(n6399), .ck(clk), .q(
        \cache_data_A[7][89] ) );
  dp_1 \cache_data_A_reg[7][90]  ( .ip(n6398), .ck(clk), .q(
        \cache_data_A[7][90] ) );
  dp_1 \cache_data_A_reg[7][91]  ( .ip(n6397), .ck(clk), .q(
        \cache_data_A[7][91] ) );
  dp_1 \cache_data_A_reg[7][92]  ( .ip(n6396), .ck(clk), .q(
        \cache_data_A[7][92] ) );
  dp_1 \cache_data_A_reg[7][93]  ( .ip(n6395), .ck(clk), .q(
        \cache_data_A[7][93] ) );
  dp_1 \cache_data_A_reg[7][94]  ( .ip(n6394), .ck(clk), .q(
        \cache_data_A[7][94] ) );
  dp_1 \cache_data_A_reg[7][95]  ( .ip(n6393), .ck(clk), .q(
        \cache_data_A[7][95] ) );
  dp_1 \cache_data_A_reg[0][124]  ( .ip(n7288), .ck(clk), .q(
        \cache_data_A[0][124] ) );
  dp_1 \cache_data_A_reg[0][125]  ( .ip(n7287), .ck(clk), .q(
        \cache_data_A[0][125] ) );
  dp_1 \cache_data_A_reg[0][126]  ( .ip(n7286), .ck(clk), .q(
        \cache_data_A[0][126] ) );
  dp_1 \cache_data_A_reg[0][127]  ( .ip(n7285), .ck(clk), .q(
        \cache_data_A[0][127] ) );
  dp_1 \cache_data_A_reg[0][96]  ( .ip(n7284), .ck(clk), .q(
        \cache_data_A[0][96] ) );
  dp_1 \cache_data_A_reg[0][97]  ( .ip(n7283), .ck(clk), .q(
        \cache_data_A[0][97] ) );
  dp_1 \cache_data_A_reg[0][98]  ( .ip(n7282), .ck(clk), .q(
        \cache_data_A[0][98] ) );
  dp_1 \cache_data_A_reg[0][99]  ( .ip(n7281), .ck(clk), .q(
        \cache_data_A[0][99] ) );
  dp_1 \cache_data_A_reg[0][100]  ( .ip(n7280), .ck(clk), .q(
        \cache_data_A[0][100] ) );
  dp_1 \cache_data_A_reg[0][101]  ( .ip(n7279), .ck(clk), .q(
        \cache_data_A[0][101] ) );
  dp_1 \cache_data_A_reg[0][102]  ( .ip(n7278), .ck(clk), .q(
        \cache_data_A[0][102] ) );
  dp_1 \cache_data_A_reg[0][103]  ( .ip(n7277), .ck(clk), .q(
        \cache_data_A[0][103] ) );
  dp_1 \cache_data_A_reg[0][104]  ( .ip(n7276), .ck(clk), .q(
        \cache_data_A[0][104] ) );
  dp_1 \cache_data_A_reg[0][105]  ( .ip(n7275), .ck(clk), .q(
        \cache_data_A[0][105] ) );
  dp_1 \cache_data_A_reg[0][106]  ( .ip(n7274), .ck(clk), .q(
        \cache_data_A[0][106] ) );
  dp_1 \cache_data_A_reg[0][107]  ( .ip(n7273), .ck(clk), .q(
        \cache_data_A[0][107] ) );
  dp_1 \cache_data_A_reg[0][108]  ( .ip(n7272), .ck(clk), .q(
        \cache_data_A[0][108] ) );
  dp_1 \cache_data_A_reg[0][109]  ( .ip(n7271), .ck(clk), .q(
        \cache_data_A[0][109] ) );
  dp_1 \cache_data_A_reg[0][110]  ( .ip(n7270), .ck(clk), .q(
        \cache_data_A[0][110] ) );
  dp_1 \cache_data_A_reg[0][111]  ( .ip(n7269), .ck(clk), .q(
        \cache_data_A[0][111] ) );
  dp_1 \cache_data_A_reg[0][112]  ( .ip(n7268), .ck(clk), .q(
        \cache_data_A[0][112] ) );
  dp_1 \cache_data_A_reg[0][113]  ( .ip(n7267), .ck(clk), .q(
        \cache_data_A[0][113] ) );
  dp_1 \cache_data_A_reg[0][114]  ( .ip(n7266), .ck(clk), .q(
        \cache_data_A[0][114] ) );
  dp_1 \cache_data_A_reg[0][115]  ( .ip(n7265), .ck(clk), .q(
        \cache_data_A[0][115] ) );
  dp_1 \cache_data_A_reg[0][116]  ( .ip(n7264), .ck(clk), .q(
        \cache_data_A[0][116] ) );
  dp_1 \cache_data_A_reg[0][117]  ( .ip(n7263), .ck(clk), .q(
        \cache_data_A[0][117] ) );
  dp_1 \cache_data_A_reg[0][118]  ( .ip(n7262), .ck(clk), .q(
        \cache_data_A[0][118] ) );
  dp_1 \cache_data_A_reg[0][119]  ( .ip(n7261), .ck(clk), .q(
        \cache_data_A[0][119] ) );
  dp_1 \cache_data_A_reg[0][120]  ( .ip(n7260), .ck(clk), .q(
        \cache_data_A[0][120] ) );
  dp_1 \cache_data_A_reg[0][121]  ( .ip(n7259), .ck(clk), .q(
        \cache_data_A[0][121] ) );
  dp_1 \cache_data_A_reg[0][122]  ( .ip(n7258), .ck(clk), .q(
        \cache_data_A[0][122] ) );
  dp_1 \cache_data_A_reg[0][123]  ( .ip(n7257), .ck(clk), .q(
        \cache_data_A[0][123] ) );
  dp_1 \cache_data_A_reg[1][96]  ( .ip(n7160), .ck(clk), .q(
        \cache_data_A[1][96] ) );
  dp_1 \cache_data_A_reg[1][97]  ( .ip(n7159), .ck(clk), .q(
        \cache_data_A[1][97] ) );
  dp_1 \cache_data_A_reg[1][98]  ( .ip(n7158), .ck(clk), .q(
        \cache_data_A[1][98] ) );
  dp_1 \cache_data_A_reg[1][99]  ( .ip(n7157), .ck(clk), .q(
        \cache_data_A[1][99] ) );
  dp_1 \cache_data_A_reg[1][100]  ( .ip(n7156), .ck(clk), .q(
        \cache_data_A[1][100] ) );
  dp_1 \cache_data_A_reg[1][101]  ( .ip(n7155), .ck(clk), .q(
        \cache_data_A[1][101] ) );
  dp_1 \cache_data_A_reg[1][102]  ( .ip(n7154), .ck(clk), .q(
        \cache_data_A[1][102] ) );
  dp_1 \cache_data_A_reg[1][103]  ( .ip(n7153), .ck(clk), .q(
        \cache_data_A[1][103] ) );
  dp_1 \cache_data_A_reg[1][104]  ( .ip(n7152), .ck(clk), .q(
        \cache_data_A[1][104] ) );
  dp_1 \cache_data_A_reg[1][105]  ( .ip(n7151), .ck(clk), .q(
        \cache_data_A[1][105] ) );
  dp_1 \cache_data_A_reg[1][106]  ( .ip(n7150), .ck(clk), .q(
        \cache_data_A[1][106] ) );
  dp_1 \cache_data_A_reg[1][107]  ( .ip(n7149), .ck(clk), .q(
        \cache_data_A[1][107] ) );
  dp_1 \cache_data_A_reg[1][108]  ( .ip(n7148), .ck(clk), .q(
        \cache_data_A[1][108] ) );
  dp_1 \cache_data_A_reg[1][109]  ( .ip(n7147), .ck(clk), .q(
        \cache_data_A[1][109] ) );
  dp_1 \cache_data_A_reg[1][110]  ( .ip(n7146), .ck(clk), .q(
        \cache_data_A[1][110] ) );
  dp_1 \cache_data_A_reg[1][111]  ( .ip(n7145), .ck(clk), .q(
        \cache_data_A[1][111] ) );
  dp_1 \cache_data_A_reg[1][112]  ( .ip(n7144), .ck(clk), .q(
        \cache_data_A[1][112] ) );
  dp_1 \cache_data_A_reg[1][113]  ( .ip(n7143), .ck(clk), .q(
        \cache_data_A[1][113] ) );
  dp_1 \cache_data_A_reg[1][114]  ( .ip(n7142), .ck(clk), .q(
        \cache_data_A[1][114] ) );
  dp_1 \cache_data_A_reg[1][115]  ( .ip(n7141), .ck(clk), .q(
        \cache_data_A[1][115] ) );
  dp_1 \cache_data_A_reg[1][116]  ( .ip(n7140), .ck(clk), .q(
        \cache_data_A[1][116] ) );
  dp_1 \cache_data_A_reg[1][117]  ( .ip(n7139), .ck(clk), .q(
        \cache_data_A[1][117] ) );
  dp_1 \cache_data_A_reg[1][118]  ( .ip(n7138), .ck(clk), .q(
        \cache_data_A[1][118] ) );
  dp_1 \cache_data_A_reg[1][119]  ( .ip(n7137), .ck(clk), .q(
        \cache_data_A[1][119] ) );
  dp_1 \cache_data_A_reg[1][120]  ( .ip(n7136), .ck(clk), .q(
        \cache_data_A[1][120] ) );
  dp_1 \cache_data_A_reg[1][121]  ( .ip(n7135), .ck(clk), .q(
        \cache_data_A[1][121] ) );
  dp_1 \cache_data_A_reg[1][122]  ( .ip(n7134), .ck(clk), .q(
        \cache_data_A[1][122] ) );
  dp_1 \cache_data_A_reg[1][123]  ( .ip(n7133), .ck(clk), .q(
        \cache_data_A[1][123] ) );
  dp_1 \cache_data_A_reg[1][124]  ( .ip(n7132), .ck(clk), .q(
        \cache_data_A[1][124] ) );
  dp_1 \cache_data_A_reg[1][125]  ( .ip(n7131), .ck(clk), .q(
        \cache_data_A[1][125] ) );
  dp_1 \cache_data_A_reg[1][126]  ( .ip(n7130), .ck(clk), .q(
        \cache_data_A[1][126] ) );
  dp_1 \cache_data_A_reg[1][127]  ( .ip(n7129), .ck(clk), .q(
        \cache_data_A[1][127] ) );
  dp_1 \cache_data_A_reg[2][96]  ( .ip(n7032), .ck(clk), .q(
        \cache_data_A[2][96] ) );
  dp_1 \cache_data_A_reg[2][97]  ( .ip(n7031), .ck(clk), .q(
        \cache_data_A[2][97] ) );
  dp_1 \cache_data_A_reg[2][98]  ( .ip(n7030), .ck(clk), .q(
        \cache_data_A[2][98] ) );
  dp_1 \cache_data_A_reg[2][99]  ( .ip(n7029), .ck(clk), .q(
        \cache_data_A[2][99] ) );
  dp_1 \cache_data_A_reg[2][100]  ( .ip(n7028), .ck(clk), .q(
        \cache_data_A[2][100] ) );
  dp_1 \cache_data_A_reg[2][101]  ( .ip(n7027), .ck(clk), .q(
        \cache_data_A[2][101] ) );
  dp_1 \cache_data_A_reg[2][102]  ( .ip(n7026), .ck(clk), .q(
        \cache_data_A[2][102] ) );
  dp_1 \cache_data_A_reg[2][103]  ( .ip(n7025), .ck(clk), .q(
        \cache_data_A[2][103] ) );
  dp_1 \cache_data_A_reg[2][104]  ( .ip(n7024), .ck(clk), .q(
        \cache_data_A[2][104] ) );
  dp_1 \cache_data_A_reg[2][105]  ( .ip(n7023), .ck(clk), .q(
        \cache_data_A[2][105] ) );
  dp_1 \cache_data_A_reg[2][106]  ( .ip(n7022), .ck(clk), .q(
        \cache_data_A[2][106] ) );
  dp_1 \cache_data_A_reg[2][107]  ( .ip(n7021), .ck(clk), .q(
        \cache_data_A[2][107] ) );
  dp_1 \cache_data_A_reg[2][108]  ( .ip(n7020), .ck(clk), .q(
        \cache_data_A[2][108] ) );
  dp_1 \cache_data_A_reg[2][109]  ( .ip(n7019), .ck(clk), .q(
        \cache_data_A[2][109] ) );
  dp_1 \cache_data_A_reg[2][110]  ( .ip(n7018), .ck(clk), .q(
        \cache_data_A[2][110] ) );
  dp_1 \cache_data_A_reg[2][111]  ( .ip(n7017), .ck(clk), .q(
        \cache_data_A[2][111] ) );
  dp_1 \cache_data_A_reg[2][112]  ( .ip(n7016), .ck(clk), .q(
        \cache_data_A[2][112] ) );
  dp_1 \cache_data_A_reg[2][113]  ( .ip(n7015), .ck(clk), .q(
        \cache_data_A[2][113] ) );
  dp_1 \cache_data_A_reg[2][114]  ( .ip(n7014), .ck(clk), .q(
        \cache_data_A[2][114] ) );
  dp_1 \cache_data_A_reg[2][115]  ( .ip(n7013), .ck(clk), .q(
        \cache_data_A[2][115] ) );
  dp_1 \cache_data_A_reg[2][116]  ( .ip(n7012), .ck(clk), .q(
        \cache_data_A[2][116] ) );
  dp_1 \cache_data_A_reg[2][117]  ( .ip(n7011), .ck(clk), .q(
        \cache_data_A[2][117] ) );
  dp_1 \cache_data_A_reg[2][118]  ( .ip(n7010), .ck(clk), .q(
        \cache_data_A[2][118] ) );
  dp_1 \cache_data_A_reg[2][119]  ( .ip(n7009), .ck(clk), .q(
        \cache_data_A[2][119] ) );
  dp_1 \cache_data_A_reg[2][120]  ( .ip(n7008), .ck(clk), .q(
        \cache_data_A[2][120] ) );
  dp_1 \cache_data_A_reg[2][121]  ( .ip(n7007), .ck(clk), .q(
        \cache_data_A[2][121] ) );
  dp_1 \cache_data_A_reg[2][122]  ( .ip(n7006), .ck(clk), .q(
        \cache_data_A[2][122] ) );
  dp_1 \cache_data_A_reg[2][123]  ( .ip(n7005), .ck(clk), .q(
        \cache_data_A[2][123] ) );
  dp_1 \cache_data_A_reg[2][124]  ( .ip(n7004), .ck(clk), .q(
        \cache_data_A[2][124] ) );
  dp_1 \cache_data_A_reg[2][125]  ( .ip(n7003), .ck(clk), .q(
        \cache_data_A[2][125] ) );
  dp_1 \cache_data_A_reg[2][126]  ( .ip(n7002), .ck(clk), .q(
        \cache_data_A[2][126] ) );
  dp_1 \cache_data_A_reg[2][127]  ( .ip(n7001), .ck(clk), .q(
        \cache_data_A[2][127] ) );
  dp_1 \cache_data_A_reg[3][96]  ( .ip(n6904), .ck(clk), .q(
        \cache_data_A[3][96] ) );
  dp_1 \cache_data_A_reg[3][97]  ( .ip(n6903), .ck(clk), .q(
        \cache_data_A[3][97] ) );
  dp_1 \cache_data_A_reg[3][98]  ( .ip(n6902), .ck(clk), .q(
        \cache_data_A[3][98] ) );
  dp_1 \cache_data_A_reg[3][99]  ( .ip(n6901), .ck(clk), .q(
        \cache_data_A[3][99] ) );
  dp_1 \cache_data_A_reg[3][100]  ( .ip(n6900), .ck(clk), .q(
        \cache_data_A[3][100] ) );
  dp_1 \cache_data_A_reg[3][101]  ( .ip(n6899), .ck(clk), .q(
        \cache_data_A[3][101] ) );
  dp_1 \cache_data_A_reg[3][102]  ( .ip(n6898), .ck(clk), .q(
        \cache_data_A[3][102] ) );
  dp_1 \cache_data_A_reg[3][103]  ( .ip(n6897), .ck(clk), .q(
        \cache_data_A[3][103] ) );
  dp_1 \cache_data_A_reg[3][104]  ( .ip(n6896), .ck(clk), .q(
        \cache_data_A[3][104] ) );
  dp_1 \cache_data_A_reg[3][105]  ( .ip(n6895), .ck(clk), .q(
        \cache_data_A[3][105] ) );
  dp_1 \cache_data_A_reg[3][106]  ( .ip(n6894), .ck(clk), .q(
        \cache_data_A[3][106] ) );
  dp_1 \cache_data_A_reg[3][107]  ( .ip(n6893), .ck(clk), .q(
        \cache_data_A[3][107] ) );
  dp_1 \cache_data_A_reg[3][108]  ( .ip(n6892), .ck(clk), .q(
        \cache_data_A[3][108] ) );
  dp_1 \cache_data_A_reg[3][109]  ( .ip(n6891), .ck(clk), .q(
        \cache_data_A[3][109] ) );
  dp_1 \cache_data_A_reg[3][110]  ( .ip(n6890), .ck(clk), .q(
        \cache_data_A[3][110] ) );
  dp_1 \cache_data_A_reg[3][111]  ( .ip(n6889), .ck(clk), .q(
        \cache_data_A[3][111] ) );
  dp_1 \cache_data_A_reg[3][112]  ( .ip(n6888), .ck(clk), .q(
        \cache_data_A[3][112] ) );
  dp_1 \cache_data_A_reg[3][113]  ( .ip(n6887), .ck(clk), .q(
        \cache_data_A[3][113] ) );
  dp_1 \cache_data_A_reg[3][114]  ( .ip(n6886), .ck(clk), .q(
        \cache_data_A[3][114] ) );
  dp_1 \cache_data_A_reg[3][115]  ( .ip(n6885), .ck(clk), .q(
        \cache_data_A[3][115] ) );
  dp_1 \cache_data_A_reg[3][116]  ( .ip(n6884), .ck(clk), .q(
        \cache_data_A[3][116] ) );
  dp_1 \cache_data_A_reg[3][117]  ( .ip(n6883), .ck(clk), .q(
        \cache_data_A[3][117] ) );
  dp_1 \cache_data_A_reg[3][118]  ( .ip(n6882), .ck(clk), .q(
        \cache_data_A[3][118] ) );
  dp_1 \cache_data_A_reg[3][119]  ( .ip(n6881), .ck(clk), .q(
        \cache_data_A[3][119] ) );
  dp_1 \cache_data_A_reg[3][120]  ( .ip(n6880), .ck(clk), .q(
        \cache_data_A[3][120] ) );
  dp_1 \cache_data_A_reg[3][121]  ( .ip(n6879), .ck(clk), .q(
        \cache_data_A[3][121] ) );
  dp_1 \cache_data_A_reg[3][122]  ( .ip(n6878), .ck(clk), .q(
        \cache_data_A[3][122] ) );
  dp_1 \cache_data_A_reg[3][123]  ( .ip(n6877), .ck(clk), .q(
        \cache_data_A[3][123] ) );
  dp_1 \cache_data_A_reg[3][124]  ( .ip(n6876), .ck(clk), .q(
        \cache_data_A[3][124] ) );
  dp_1 \cache_data_A_reg[3][125]  ( .ip(n6875), .ck(clk), .q(
        \cache_data_A[3][125] ) );
  dp_1 \cache_data_A_reg[3][126]  ( .ip(n6874), .ck(clk), .q(
        \cache_data_A[3][126] ) );
  dp_1 \cache_data_A_reg[3][127]  ( .ip(n6873), .ck(clk), .q(
        \cache_data_A[3][127] ) );
  dp_1 \cache_data_A_reg[4][107]  ( .ip(n6776), .ck(clk), .q(
        \cache_data_A[4][107] ) );
  dp_1 \cache_data_A_reg[4][108]  ( .ip(n6775), .ck(clk), .q(
        \cache_data_A[4][108] ) );
  dp_1 \cache_data_A_reg[4][109]  ( .ip(n6774), .ck(clk), .q(
        \cache_data_A[4][109] ) );
  dp_1 \cache_data_A_reg[4][110]  ( .ip(n6773), .ck(clk), .q(
        \cache_data_A[4][110] ) );
  dp_1 \cache_data_A_reg[4][111]  ( .ip(n6772), .ck(clk), .q(
        \cache_data_A[4][111] ) );
  dp_1 \cache_data_A_reg[4][112]  ( .ip(n6771), .ck(clk), .q(
        \cache_data_A[4][112] ) );
  dp_1 \cache_data_A_reg[4][113]  ( .ip(n6770), .ck(clk), .q(
        \cache_data_A[4][113] ) );
  dp_1 \cache_data_A_reg[4][114]  ( .ip(n6769), .ck(clk), .q(
        \cache_data_A[4][114] ) );
  dp_1 \cache_data_A_reg[4][115]  ( .ip(n6768), .ck(clk), .q(
        \cache_data_A[4][115] ) );
  dp_1 \cache_data_A_reg[4][116]  ( .ip(n6767), .ck(clk), .q(
        \cache_data_A[4][116] ) );
  dp_1 \cache_data_A_reg[4][117]  ( .ip(n6766), .ck(clk), .q(
        \cache_data_A[4][117] ) );
  dp_1 \cache_data_A_reg[4][118]  ( .ip(n6765), .ck(clk), .q(
        \cache_data_A[4][118] ) );
  dp_1 \cache_data_A_reg[4][119]  ( .ip(n6764), .ck(clk), .q(
        \cache_data_A[4][119] ) );
  dp_1 \cache_data_A_reg[4][120]  ( .ip(n6763), .ck(clk), .q(
        \cache_data_A[4][120] ) );
  dp_1 \cache_data_A_reg[4][121]  ( .ip(n6762), .ck(clk), .q(
        \cache_data_A[4][121] ) );
  dp_1 \cache_data_A_reg[4][122]  ( .ip(n6761), .ck(clk), .q(
        \cache_data_A[4][122] ) );
  dp_1 \cache_data_A_reg[4][123]  ( .ip(n6760), .ck(clk), .q(
        \cache_data_A[4][123] ) );
  dp_1 \cache_data_A_reg[4][124]  ( .ip(n6759), .ck(clk), .q(
        \cache_data_A[4][124] ) );
  dp_1 \cache_data_A_reg[4][125]  ( .ip(n6758), .ck(clk), .q(
        \cache_data_A[4][125] ) );
  dp_1 \cache_data_A_reg[4][126]  ( .ip(n6757), .ck(clk), .q(
        \cache_data_A[4][126] ) );
  dp_1 \cache_data_A_reg[4][127]  ( .ip(n6756), .ck(clk), .q(
        \cache_data_A[4][127] ) );
  dp_1 \cache_data_A_reg[4][96]  ( .ip(n6755), .ck(clk), .q(
        \cache_data_A[4][96] ) );
  dp_1 \cache_data_A_reg[4][97]  ( .ip(n6754), .ck(clk), .q(
        \cache_data_A[4][97] ) );
  dp_1 \cache_data_A_reg[4][98]  ( .ip(n6753), .ck(clk), .q(
        \cache_data_A[4][98] ) );
  dp_1 \cache_data_A_reg[4][99]  ( .ip(n6752), .ck(clk), .q(
        \cache_data_A[4][99] ) );
  dp_1 \cache_data_A_reg[4][100]  ( .ip(n6751), .ck(clk), .q(
        \cache_data_A[4][100] ) );
  dp_1 \cache_data_A_reg[4][101]  ( .ip(n6750), .ck(clk), .q(
        \cache_data_A[4][101] ) );
  dp_1 \cache_data_A_reg[4][102]  ( .ip(n6749), .ck(clk), .q(
        \cache_data_A[4][102] ) );
  dp_1 \cache_data_A_reg[4][103]  ( .ip(n6748), .ck(clk), .q(
        \cache_data_A[4][103] ) );
  dp_1 \cache_data_A_reg[4][104]  ( .ip(n6747), .ck(clk), .q(
        \cache_data_A[4][104] ) );
  dp_1 \cache_data_A_reg[4][105]  ( .ip(n6746), .ck(clk), .q(
        \cache_data_A[4][105] ) );
  dp_1 \cache_data_A_reg[4][106]  ( .ip(n6745), .ck(clk), .q(
        \cache_data_A[4][106] ) );
  dp_1 \cache_data_A_reg[5][96]  ( .ip(n6648), .ck(clk), .q(
        \cache_data_A[5][96] ) );
  dp_1 \cache_data_A_reg[5][97]  ( .ip(n6647), .ck(clk), .q(
        \cache_data_A[5][97] ) );
  dp_1 \cache_data_A_reg[5][98]  ( .ip(n6646), .ck(clk), .q(
        \cache_data_A[5][98] ) );
  dp_1 \cache_data_A_reg[5][99]  ( .ip(n6645), .ck(clk), .q(
        \cache_data_A[5][99] ) );
  dp_1 \cache_data_A_reg[5][100]  ( .ip(n6644), .ck(clk), .q(
        \cache_data_A[5][100] ) );
  dp_1 \cache_data_A_reg[5][101]  ( .ip(n6643), .ck(clk), .q(
        \cache_data_A[5][101] ) );
  dp_1 \cache_data_A_reg[5][102]  ( .ip(n6642), .ck(clk), .q(
        \cache_data_A[5][102] ) );
  dp_1 \cache_data_A_reg[5][103]  ( .ip(n6641), .ck(clk), .q(
        \cache_data_A[5][103] ) );
  dp_1 \cache_data_A_reg[5][104]  ( .ip(n6640), .ck(clk), .q(
        \cache_data_A[5][104] ) );
  dp_1 \cache_data_A_reg[5][105]  ( .ip(n6639), .ck(clk), .q(
        \cache_data_A[5][105] ) );
  dp_1 \cache_data_A_reg[5][106]  ( .ip(n6638), .ck(clk), .q(
        \cache_data_A[5][106] ) );
  dp_1 \cache_data_A_reg[5][107]  ( .ip(n6637), .ck(clk), .q(
        \cache_data_A[5][107] ) );
  dp_1 \cache_data_A_reg[5][108]  ( .ip(n6636), .ck(clk), .q(
        \cache_data_A[5][108] ) );
  dp_1 \cache_data_A_reg[5][109]  ( .ip(n6635), .ck(clk), .q(
        \cache_data_A[5][109] ) );
  dp_1 \cache_data_A_reg[5][110]  ( .ip(n6634), .ck(clk), .q(
        \cache_data_A[5][110] ) );
  dp_1 \cache_data_A_reg[5][111]  ( .ip(n6633), .ck(clk), .q(
        \cache_data_A[5][111] ) );
  dp_1 \cache_data_A_reg[5][112]  ( .ip(n6632), .ck(clk), .q(
        \cache_data_A[5][112] ) );
  dp_1 \cache_data_A_reg[5][113]  ( .ip(n6631), .ck(clk), .q(
        \cache_data_A[5][113] ) );
  dp_1 \cache_data_A_reg[5][114]  ( .ip(n6630), .ck(clk), .q(
        \cache_data_A[5][114] ) );
  dp_1 \cache_data_A_reg[5][115]  ( .ip(n6629), .ck(clk), .q(
        \cache_data_A[5][115] ) );
  dp_1 \cache_data_A_reg[5][116]  ( .ip(n6628), .ck(clk), .q(
        \cache_data_A[5][116] ) );
  dp_1 \cache_data_A_reg[5][117]  ( .ip(n6627), .ck(clk), .q(
        \cache_data_A[5][117] ) );
  dp_1 \cache_data_A_reg[5][118]  ( .ip(n6626), .ck(clk), .q(
        \cache_data_A[5][118] ) );
  dp_1 \cache_data_A_reg[5][119]  ( .ip(n6625), .ck(clk), .q(
        \cache_data_A[5][119] ) );
  dp_1 \cache_data_A_reg[5][120]  ( .ip(n6624), .ck(clk), .q(
        \cache_data_A[5][120] ) );
  dp_1 \cache_data_A_reg[5][121]  ( .ip(n6623), .ck(clk), .q(
        \cache_data_A[5][121] ) );
  dp_1 \cache_data_A_reg[5][122]  ( .ip(n6622), .ck(clk), .q(
        \cache_data_A[5][122] ) );
  dp_1 \cache_data_A_reg[5][123]  ( .ip(n6621), .ck(clk), .q(
        \cache_data_A[5][123] ) );
  dp_1 \cache_data_A_reg[5][124]  ( .ip(n6620), .ck(clk), .q(
        \cache_data_A[5][124] ) );
  dp_1 \cache_data_A_reg[5][125]  ( .ip(n6619), .ck(clk), .q(
        \cache_data_A[5][125] ) );
  dp_1 \cache_data_A_reg[5][126]  ( .ip(n6618), .ck(clk), .q(
        \cache_data_A[5][126] ) );
  dp_1 \cache_data_A_reg[5][127]  ( .ip(n6617), .ck(clk), .q(
        \cache_data_A[5][127] ) );
  dp_1 \cache_data_A_reg[6][96]  ( .ip(n6520), .ck(clk), .q(
        \cache_data_A[6][96] ) );
  dp_1 \cache_data_A_reg[6][97]  ( .ip(n6519), .ck(clk), .q(
        \cache_data_A[6][97] ) );
  dp_1 \cache_data_A_reg[6][98]  ( .ip(n6518), .ck(clk), .q(
        \cache_data_A[6][98] ) );
  dp_1 \cache_data_A_reg[6][99]  ( .ip(n6517), .ck(clk), .q(
        \cache_data_A[6][99] ) );
  dp_1 \cache_data_A_reg[6][100]  ( .ip(n6516), .ck(clk), .q(
        \cache_data_A[6][100] ) );
  dp_1 \cache_data_A_reg[6][101]  ( .ip(n6515), .ck(clk), .q(
        \cache_data_A[6][101] ) );
  dp_1 \cache_data_A_reg[6][102]  ( .ip(n6514), .ck(clk), .q(
        \cache_data_A[6][102] ) );
  dp_1 \cache_data_A_reg[6][103]  ( .ip(n6513), .ck(clk), .q(
        \cache_data_A[6][103] ) );
  dp_1 \cache_data_A_reg[6][104]  ( .ip(n6512), .ck(clk), .q(
        \cache_data_A[6][104] ) );
  dp_1 \cache_data_A_reg[6][105]  ( .ip(n6511), .ck(clk), .q(
        \cache_data_A[6][105] ) );
  dp_1 \cache_data_A_reg[6][106]  ( .ip(n6510), .ck(clk), .q(
        \cache_data_A[6][106] ) );
  dp_1 \cache_data_A_reg[6][107]  ( .ip(n6509), .ck(clk), .q(
        \cache_data_A[6][107] ) );
  dp_1 \cache_data_A_reg[6][108]  ( .ip(n6508), .ck(clk), .q(
        \cache_data_A[6][108] ) );
  dp_1 \cache_data_A_reg[6][109]  ( .ip(n6507), .ck(clk), .q(
        \cache_data_A[6][109] ) );
  dp_1 \cache_data_A_reg[6][110]  ( .ip(n6506), .ck(clk), .q(
        \cache_data_A[6][110] ) );
  dp_1 \cache_data_A_reg[6][111]  ( .ip(n6505), .ck(clk), .q(
        \cache_data_A[6][111] ) );
  dp_1 \cache_data_A_reg[6][112]  ( .ip(n6504), .ck(clk), .q(
        \cache_data_A[6][112] ) );
  dp_1 \cache_data_A_reg[6][113]  ( .ip(n6503), .ck(clk), .q(
        \cache_data_A[6][113] ) );
  dp_1 \cache_data_A_reg[6][114]  ( .ip(n6502), .ck(clk), .q(
        \cache_data_A[6][114] ) );
  dp_1 \cache_data_A_reg[6][115]  ( .ip(n6501), .ck(clk), .q(
        \cache_data_A[6][115] ) );
  dp_1 \cache_data_A_reg[6][116]  ( .ip(n6500), .ck(clk), .q(
        \cache_data_A[6][116] ) );
  dp_1 \cache_data_A_reg[6][117]  ( .ip(n6499), .ck(clk), .q(
        \cache_data_A[6][117] ) );
  dp_1 \cache_data_A_reg[6][118]  ( .ip(n6498), .ck(clk), .q(
        \cache_data_A[6][118] ) );
  dp_1 \cache_data_A_reg[6][119]  ( .ip(n6497), .ck(clk), .q(
        \cache_data_A[6][119] ) );
  dp_1 \cache_data_A_reg[6][120]  ( .ip(n6496), .ck(clk), .q(
        \cache_data_A[6][120] ) );
  dp_1 \cache_data_A_reg[6][121]  ( .ip(n6495), .ck(clk), .q(
        \cache_data_A[6][121] ) );
  dp_1 \cache_data_A_reg[6][122]  ( .ip(n6494), .ck(clk), .q(
        \cache_data_A[6][122] ) );
  dp_1 \cache_data_A_reg[6][123]  ( .ip(n6493), .ck(clk), .q(
        \cache_data_A[6][123] ) );
  dp_1 \cache_data_A_reg[6][124]  ( .ip(n6492), .ck(clk), .q(
        \cache_data_A[6][124] ) );
  dp_1 \cache_data_A_reg[6][125]  ( .ip(n6491), .ck(clk), .q(
        \cache_data_A[6][125] ) );
  dp_1 \cache_data_A_reg[6][126]  ( .ip(n6490), .ck(clk), .q(
        \cache_data_A[6][126] ) );
  dp_1 \cache_data_A_reg[6][127]  ( .ip(n6489), .ck(clk), .q(
        \cache_data_A[6][127] ) );
  dp_1 \cache_data_A_reg[7][119]  ( .ip(n6392), .ck(clk), .q(
        \cache_data_A[7][119] ) );
  dp_1 \data_wr_mem_reg[23]  ( .ip(n5265), .ck(clk), .q(data_wr_mem[23]) );
  dp_1 \cache_data_A_reg[7][120]  ( .ip(n6391), .ck(clk), .q(
        \cache_data_A[7][120] ) );
  dp_1 \data_wr_mem_reg[24]  ( .ip(n5264), .ck(clk), .q(data_wr_mem[24]) );
  dp_1 \cache_data_A_reg[7][121]  ( .ip(n6390), .ck(clk), .q(
        \cache_data_A[7][121] ) );
  dp_1 \data_wr_mem_reg[25]  ( .ip(n5263), .ck(clk), .q(data_wr_mem[25]) );
  dp_1 \cache_data_A_reg[7][122]  ( .ip(n6389), .ck(clk), .q(
        \cache_data_A[7][122] ) );
  dp_1 \data_wr_mem_reg[26]  ( .ip(n5262), .ck(clk), .q(data_wr_mem[26]) );
  dp_1 \cache_data_A_reg[7][123]  ( .ip(n6388), .ck(clk), .q(
        \cache_data_A[7][123] ) );
  dp_1 \data_wr_mem_reg[27]  ( .ip(n5261), .ck(clk), .q(data_wr_mem[27]) );
  dp_1 \cache_data_A_reg[7][124]  ( .ip(n6387), .ck(clk), .q(
        \cache_data_A[7][124] ) );
  dp_1 \data_wr_mem_reg[28]  ( .ip(n5260), .ck(clk), .q(data_wr_mem[28]) );
  dp_1 \cache_data_A_reg[7][125]  ( .ip(n6386), .ck(clk), .q(
        \cache_data_A[7][125] ) );
  dp_1 \data_wr_mem_reg[29]  ( .ip(n5259), .ck(clk), .q(data_wr_mem[29]) );
  dp_1 \cache_data_A_reg[7][126]  ( .ip(n6385), .ck(clk), .q(
        \cache_data_A[7][126] ) );
  dp_1 \data_wr_mem_reg[30]  ( .ip(n5258), .ck(clk), .q(data_wr_mem[30]) );
  dp_1 \cache_data_A_reg[7][127]  ( .ip(n6384), .ck(clk), .q(
        \cache_data_A[7][127] ) );
  dp_1 \data_wr_mem_reg[31]  ( .ip(n5257), .ck(clk), .q(data_wr_mem[31]) );
  dp_1 \cache_data_A_reg[7][96]  ( .ip(n6383), .ck(clk), .q(
        \cache_data_A[7][96] ) );
  dp_1 \data_wr_mem_reg[0]  ( .ip(n5288), .ck(clk), .q(data_wr_mem[0]) );
  dp_1 \cache_data_A_reg[7][97]  ( .ip(n6382), .ck(clk), .q(
        \cache_data_A[7][97] ) );
  dp_1 \data_wr_mem_reg[1]  ( .ip(n5287), .ck(clk), .q(data_wr_mem[1]) );
  dp_1 \cache_data_A_reg[7][98]  ( .ip(n6381), .ck(clk), .q(
        \cache_data_A[7][98] ) );
  dp_1 \data_wr_mem_reg[2]  ( .ip(n5286), .ck(clk), .q(data_wr_mem[2]) );
  dp_1 \cache_data_A_reg[7][99]  ( .ip(n6380), .ck(clk), .q(
        \cache_data_A[7][99] ) );
  dp_1 \data_wr_mem_reg[3]  ( .ip(n5285), .ck(clk), .q(data_wr_mem[3]) );
  dp_1 \cache_data_A_reg[7][100]  ( .ip(n6379), .ck(clk), .q(
        \cache_data_A[7][100] ) );
  dp_1 \data_wr_mem_reg[4]  ( .ip(n5284), .ck(clk), .q(data_wr_mem[4]) );
  dp_1 \cache_data_A_reg[7][101]  ( .ip(n6378), .ck(clk), .q(
        \cache_data_A[7][101] ) );
  dp_1 \data_wr_mem_reg[5]  ( .ip(n5283), .ck(clk), .q(data_wr_mem[5]) );
  dp_1 \cache_data_A_reg[7][102]  ( .ip(n6377), .ck(clk), .q(
        \cache_data_A[7][102] ) );
  dp_1 \data_wr_mem_reg[6]  ( .ip(n5282), .ck(clk), .q(data_wr_mem[6]) );
  dp_1 \cache_data_A_reg[7][103]  ( .ip(n6376), .ck(clk), .q(
        \cache_data_A[7][103] ) );
  dp_1 \data_wr_mem_reg[7]  ( .ip(n5281), .ck(clk), .q(data_wr_mem[7]) );
  dp_1 \cache_data_A_reg[7][104]  ( .ip(n6375), .ck(clk), .q(
        \cache_data_A[7][104] ) );
  dp_1 \data_wr_mem_reg[8]  ( .ip(n5280), .ck(clk), .q(data_wr_mem[8]) );
  dp_1 \cache_data_A_reg[7][105]  ( .ip(n6374), .ck(clk), .q(
        \cache_data_A[7][105] ) );
  dp_1 \data_wr_mem_reg[9]  ( .ip(n5279), .ck(clk), .q(data_wr_mem[9]) );
  dp_1 \cache_data_A_reg[7][106]  ( .ip(n6373), .ck(clk), .q(
        \cache_data_A[7][106] ) );
  dp_1 \data_wr_mem_reg[10]  ( .ip(n5278), .ck(clk), .q(data_wr_mem[10]) );
  dp_1 \cache_data_A_reg[7][107]  ( .ip(n6372), .ck(clk), .q(
        \cache_data_A[7][107] ) );
  dp_1 \data_wr_mem_reg[11]  ( .ip(n5277), .ck(clk), .q(data_wr_mem[11]) );
  dp_1 \cache_data_A_reg[7][108]  ( .ip(n6371), .ck(clk), .q(
        \cache_data_A[7][108] ) );
  dp_1 \data_wr_mem_reg[12]  ( .ip(n5276), .ck(clk), .q(data_wr_mem[12]) );
  dp_1 \cache_data_A_reg[7][109]  ( .ip(n6370), .ck(clk), .q(
        \cache_data_A[7][109] ) );
  dp_1 \data_wr_mem_reg[13]  ( .ip(n5275), .ck(clk), .q(data_wr_mem[13]) );
  dp_1 \cache_data_A_reg[7][110]  ( .ip(n6369), .ck(clk), .q(
        \cache_data_A[7][110] ) );
  dp_1 \data_wr_mem_reg[14]  ( .ip(n5274), .ck(clk), .q(data_wr_mem[14]) );
  dp_1 \cache_data_A_reg[7][111]  ( .ip(n6368), .ck(clk), .q(
        \cache_data_A[7][111] ) );
  dp_1 \data_wr_mem_reg[15]  ( .ip(n5273), .ck(clk), .q(data_wr_mem[15]) );
  dp_1 \cache_data_A_reg[7][112]  ( .ip(n6367), .ck(clk), .q(
        \cache_data_A[7][112] ) );
  dp_1 \data_wr_mem_reg[16]  ( .ip(n5272), .ck(clk), .q(data_wr_mem[16]) );
  dp_1 \cache_data_A_reg[7][113]  ( .ip(n6366), .ck(clk), .q(
        \cache_data_A[7][113] ) );
  dp_1 \data_wr_mem_reg[17]  ( .ip(n5271), .ck(clk), .q(data_wr_mem[17]) );
  dp_1 \cache_data_A_reg[7][114]  ( .ip(n6365), .ck(clk), .q(
        \cache_data_A[7][114] ) );
  dp_1 \data_wr_mem_reg[18]  ( .ip(n5270), .ck(clk), .q(data_wr_mem[18]) );
  dp_1 \cache_data_A_reg[7][115]  ( .ip(n6364), .ck(clk), .q(
        \cache_data_A[7][115] ) );
  dp_1 \data_wr_mem_reg[19]  ( .ip(n5269), .ck(clk), .q(data_wr_mem[19]) );
  dp_1 \cache_data_A_reg[7][116]  ( .ip(n6363), .ck(clk), .q(
        \cache_data_A[7][116] ) );
  dp_1 \data_wr_mem_reg[20]  ( .ip(n5268), .ck(clk), .q(data_wr_mem[20]) );
  dp_1 \cache_data_A_reg[7][117]  ( .ip(n6362), .ck(clk), .q(
        \cache_data_A[7][117] ) );
  dp_1 \data_wr_mem_reg[21]  ( .ip(n5267), .ck(clk), .q(data_wr_mem[21]) );
  dp_1 \cache_data_A_reg[7][118]  ( .ip(n6361), .ck(clk), .q(
        \cache_data_A[7][118] ) );
  dp_1 \data_wr_mem_reg[22]  ( .ip(n5266), .ck(clk), .q(data_wr_mem[22]) );
  dp_1 \data_rd_reg[0]  ( .ip(n5320), .ck(clk), .q(N4204) );
  dp_1 \data_rd_reg[1]  ( .ip(n5319), .ck(clk), .q(N4201) );
  dp_1 \data_rd_reg[2]  ( .ip(n5318), .ck(clk), .q(N4198) );
  dp_1 \data_rd_reg[3]  ( .ip(n5317), .ck(clk), .q(N4195) );
  dp_1 \data_rd_reg[4]  ( .ip(n5316), .ck(clk), .q(N4192) );
  dp_1 \data_rd_reg[5]  ( .ip(n5315), .ck(clk), .q(N4189) );
  dp_1 \data_rd_reg[6]  ( .ip(n5314), .ck(clk), .q(N4186) );
  dp_1 \data_rd_reg[7]  ( .ip(n5313), .ck(clk), .q(N4183) );
  dp_1 \data_rd_reg[8]  ( .ip(n5312), .ck(clk), .q(N4180) );
  dp_1 \data_rd_reg[9]  ( .ip(n5311), .ck(clk), .q(N4177) );
  dp_1 \data_rd_reg[10]  ( .ip(n5310), .ck(clk), .q(N4174) );
  dp_1 \data_rd_reg[11]  ( .ip(n5309), .ck(clk), .q(N4171) );
  dp_1 \data_rd_reg[12]  ( .ip(n5308), .ck(clk), .q(N4168) );
  dp_1 \data_rd_reg[13]  ( .ip(n5307), .ck(clk), .q(N4165) );
  dp_1 \data_rd_reg[14]  ( .ip(n5306), .ck(clk), .q(N4162) );
  dp_1 \data_rd_reg[15]  ( .ip(n5305), .ck(clk), .q(N4159) );
  dp_1 \data_rd_reg[16]  ( .ip(n5304), .ck(clk), .q(N4156) );
  dp_1 \data_rd_reg[17]  ( .ip(n5303), .ck(clk), .q(N4153) );
  dp_1 \data_rd_reg[18]  ( .ip(n5302), .ck(clk), .q(N4150) );
  dp_1 \data_rd_reg[19]  ( .ip(n5301), .ck(clk), .q(N4147) );
  dp_1 \data_rd_reg[20]  ( .ip(n5300), .ck(clk), .q(N4144) );
  dp_1 \data_rd_reg[21]  ( .ip(n5299), .ck(clk), .q(N4141) );
  dp_1 \data_rd_reg[22]  ( .ip(n5298), .ck(clk), .q(N4138) );
  dp_1 \data_rd_reg[23]  ( .ip(n5297), .ck(clk), .q(N4135) );
  dp_1 \data_rd_reg[24]  ( .ip(n5296), .ck(clk), .q(N4132) );
  dp_1 \data_rd_reg[25]  ( .ip(n5295), .ck(clk), .q(N4129) );
  dp_1 \data_rd_reg[26]  ( .ip(n5294), .ck(clk), .q(N4126) );
  dp_1 \data_rd_reg[27]  ( .ip(n5293), .ck(clk), .q(N4123) );
  dp_1 \data_rd_reg[28]  ( .ip(n5292), .ck(clk), .q(N4120) );
  dp_1 \data_rd_reg[29]  ( .ip(n5291), .ck(clk), .q(N4117) );
  dp_1 \data_rd_reg[30]  ( .ip(n5290), .ck(clk), .q(N4114) );
  dp_1 \data_rd_reg[31]  ( .ip(n5289), .ck(clk), .q(N4111) );
  invzp_1 \data_rd_tri[0]  ( .ip(n63), .c(N4205), .op(data_rd[0]) );
  invzp_1 \data_rd_tri[1]  ( .ip(n61), .c(N4202), .op(data_rd[1]) );
  invzp_1 \data_rd_tri[2]  ( .ip(n59), .c(N4199), .op(data_rd[2]) );
  invzp_1 \data_rd_tri[3]  ( .ip(n57), .c(N4196), .op(data_rd[3]) );
  invzp_1 \data_rd_tri[4]  ( .ip(n55), .c(N4193), .op(data_rd[4]) );
  invzp_1 \data_rd_tri[5]  ( .ip(n53), .c(N4190), .op(data_rd[5]) );
  invzp_1 \data_rd_tri[6]  ( .ip(n51), .c(N4187), .op(data_rd[6]) );
  invzp_1 \data_rd_tri[7]  ( .ip(n49), .c(N4184), .op(data_rd[7]) );
  invzp_1 \data_rd_tri[8]  ( .ip(n47), .c(N4181), .op(data_rd[8]) );
  invzp_1 \data_rd_tri[9]  ( .ip(n45), .c(N4178), .op(data_rd[9]) );
  invzp_1 \data_rd_tri[10]  ( .ip(n43), .c(N4175), .op(data_rd[10]) );
  invzp_1 \data_rd_tri[11]  ( .ip(n41), .c(N4172), .op(data_rd[11]) );
  invzp_1 \data_rd_tri[12]  ( .ip(n39), .c(N4169), .op(data_rd[12]) );
  invzp_1 \data_rd_tri[13]  ( .ip(n37), .c(N4166), .op(data_rd[13]) );
  invzp_1 \data_rd_tri[14]  ( .ip(n35), .c(N4163), .op(data_rd[14]) );
  invzp_1 \data_rd_tri[15]  ( .ip(n33), .c(N4160), .op(data_rd[15]) );
  invzp_1 \data_rd_tri[16]  ( .ip(n31), .c(N4157), .op(data_rd[16]) );
  invzp_1 \data_rd_tri[17]  ( .ip(n29), .c(N4154), .op(data_rd[17]) );
  invzp_1 \data_rd_tri[18]  ( .ip(n27), .c(N4151), .op(data_rd[18]) );
  invzp_1 \data_rd_tri[19]  ( .ip(n25), .c(N4148), .op(data_rd[19]) );
  invzp_1 \data_rd_tri[20]  ( .ip(n23), .c(N4145), .op(data_rd[20]) );
  invzp_1 \data_rd_tri[21]  ( .ip(n21), .c(N4142), .op(data_rd[21]) );
  invzp_1 \data_rd_tri[22]  ( .ip(n19), .c(N4139), .op(data_rd[22]) );
  invzp_1 \data_rd_tri[23]  ( .ip(n17), .c(N4136), .op(data_rd[23]) );
  invzp_1 \data_rd_tri[24]  ( .ip(n15), .c(N4133), .op(data_rd[24]) );
  invzp_1 \data_rd_tri[25]  ( .ip(n13), .c(N4130), .op(data_rd[25]) );
  invzp_1 \data_rd_tri[26]  ( .ip(n11), .c(N4127), .op(data_rd[26]) );
  invzp_1 \data_rd_tri[27]  ( .ip(n9), .c(N4124), .op(data_rd[27]) );
  invzp_1 \data_rd_tri[28]  ( .ip(n7), .c(N4121), .op(data_rd[28]) );
  invzp_1 \data_rd_tri[29]  ( .ip(n5), .c(N4118), .op(data_rd[29]) );
  invzp_1 \data_rd_tri[30]  ( .ip(n3), .c(N4115), .op(data_rd[30]) );
  invzp_1 \data_rd_tri[31]  ( .ip(n1), .c(N4112), .op(data_rd[31]) );
  invzp_1 \addr_resp_tri[0]  ( .ip(n127), .c(N4301), .op(addr_resp[0]) );
  invzp_1 \addr_resp_tri[1]  ( .ip(n125), .c(N4298), .op(addr_resp[1]) );
  invzp_1 \addr_resp_tri[3]  ( .ip(n121), .c(N4292), .op(addr_resp[3]) );
  invzp_1 \addr_resp_tri[2]  ( .ip(n123), .c(N4295), .op(addr_resp[2]) );
  invzp_1 \addr_resp_tri[25]  ( .ip(n77), .c(N4226), .op(addr_resp[25]) );
  invzp_1 \addr_resp_tri[15]  ( .ip(n97), .c(N4256), .op(addr_resp[15]) );
  invzp_1 \addr_resp_tri[21]  ( .ip(n85), .c(N4238), .op(addr_resp[21]) );
  invzp_1 \addr_resp_tri[24]  ( .ip(n79), .c(N4229), .op(addr_resp[24]) );
  invzp_1 \addr_resp_tri[28]  ( .ip(n71), .c(N4217), .op(addr_resp[28]) );
  invzp_1 \addr_resp_tri[26]  ( .ip(n75), .c(N4223), .op(addr_resp[26]) );
  invzp_1 \addr_resp_tri[14]  ( .ip(n99), .c(N4259), .op(addr_resp[14]) );
  invzp_1 \addr_resp_tri[19]  ( .ip(n89), .c(N4244), .op(addr_resp[19]) );
  invzp_1 \addr_resp_tri[30]  ( .ip(n67), .c(N4211), .op(addr_resp[30]) );
  invzp_1 \addr_resp_tri[10]  ( .ip(n107), .c(N4271), .op(addr_resp[10]) );
  invzp_1 \addr_resp_tri[17]  ( .ip(n93), .c(N4250), .op(addr_resp[17]) );
  invzp_1 \addr_resp_tri[16]  ( .ip(n95), .c(N4253), .op(addr_resp[16]) );
  invzp_1 \addr_resp_tri[18]  ( .ip(n91), .c(N4247), .op(addr_resp[18]) );
  invzp_1 \addr_resp_tri[20]  ( .ip(n87), .c(N4241), .op(addr_resp[20]) );
  invzp_1 \addr_resp_tri[29]  ( .ip(n69), .c(N4214), .op(addr_resp[29]) );
  invzp_1 \addr_resp_tri[13]  ( .ip(n101), .c(N4262), .op(addr_resp[13]) );
  invzp_1 \addr_resp_tri[22]  ( .ip(n83), .c(N4235), .op(addr_resp[22]) );
  invzp_1 \addr_resp_tri[31]  ( .ip(n65), .c(N4208), .op(addr_resp[31]) );
  invzp_1 \addr_resp_tri[8]  ( .ip(n111), .c(N4277), .op(addr_resp[8]) );
  invzp_1 \addr_resp_tri[9]  ( .ip(n109), .c(N4274), .op(addr_resp[9]) );
  invzp_1 \addr_resp_tri[12]  ( .ip(n103), .c(N4265), .op(addr_resp[12]) );
  invzp_1 \addr_resp_tri[23]  ( .ip(n81), .c(N4232), .op(addr_resp[23]) );
  invzp_1 \addr_resp_tri[7]  ( .ip(n113), .c(N4280), .op(addr_resp[7]) );
  invzp_1 \addr_resp_tri[11]  ( .ip(n105), .c(N4268), .op(addr_resp[11]) );
  invzp_1 \addr_resp_tri[27]  ( .ip(n73), .c(N4220), .op(addr_resp[27]) );
  invzp_1 \addr_resp_tri[4]  ( .ip(n119), .c(N4289), .op(addr_resp[4]) );
  invzp_1 \addr_resp_tri[6]  ( .ip(n115), .c(N4283), .op(addr_resp[6]) );
  invzp_1 \addr_resp_tri[5]  ( .ip(n117), .c(N4286), .op(addr_resp[5]) );
  drp_1 \cache_miss_count_reg[0]  ( .ip(n5189), .ck(clk), .rb(n7947), .q(
        cache_miss_count[0]) );
  drp_1 \cache_hit_count_reg[1]  ( .ip(n5157), .ck(clk), .rb(n7945), .q(
        cache_hit_count[1]) );
  drp_1 \cache_hit_count_reg[0]  ( .ip(n5156), .ck(clk), .rb(n7944), .q(
        cache_hit_count[0]) );
  drp_1 \state_reg[2]  ( .ip(next_state[2]), .ck(clk), .rb(n7945), .q(state[2]) );
  drp_1 \cache_miss_count_reg[1]  ( .ip(n5190), .ck(clk), .rb(n7945), .q(
        cache_miss_count[1]) );
  drp_1 \state_reg[1]  ( .ip(next_state[1]), .ck(clk), .rb(n7949), .q(state[1]) );
  drp_1 \cache_miss_count_reg[2]  ( .ip(n5191), .ck(clk), .rb(n7947), .q(
        cache_miss_count[2]) );
  drp_1 \cache_hit_count_reg[3]  ( .ip(n5159), .ck(clk), .rb(n7945), .q(
        cache_hit_count[3]) );
  drp_1 \cache_hit_count_reg[2]  ( .ip(n5158), .ck(clk), .rb(n7947), .q(
        cache_hit_count[2]) );
  drp_1 \state_reg[4]  ( .ip(n13294), .ck(clk), .rb(n7950), .q(state[4]) );
  drp_1 rdy_reg ( .ip(n13294), .ck(clk), .rb(n7947), .q(rdy) );
  drp_1 \cache_miss_count_reg[3]  ( .ip(n5192), .ck(clk), .rb(n7947), .q(
        cache_miss_count[3]) );
  drp_1 \cache_miss_count_reg[4]  ( .ip(n5193), .ck(clk), .rb(n7943), .q(
        cache_miss_count[4]) );
  drp_1 \cache_hit_count_reg[5]  ( .ip(n5161), .ck(clk), .rb(n7948), .q(
        cache_hit_count[5]) );
  drp_1 \cache_hit_count_reg[4]  ( .ip(n5160), .ck(clk), .rb(n7947), .q(
        cache_hit_count[4]) );
  drp_1 \state_reg[3]  ( .ip(n13295), .ck(clk), .rb(n7950), .q(state[3]) );
  drp_1 \cache_miss_count_reg[5]  ( .ip(n5194), .ck(clk), .rb(n7945), .q(
        cache_miss_count[5]) );
  drp_1 \cache_hit_count_reg[7]  ( .ip(n5163), .ck(clk), .rb(n7949), .q(
        cache_hit_count[7]) );
  drp_1 \cache_miss_count_reg[6]  ( .ip(n5195), .ck(clk), .rb(n7950), .q(
        cache_miss_count[6]) );
  drp_1 \cache_hit_count_reg[6]  ( .ip(n5162), .ck(clk), .rb(n7950), .q(
        cache_hit_count[6]) );
  drp_1 \cache_miss_count_reg[7]  ( .ip(n5196), .ck(clk), .rb(n7947), .q(
        cache_miss_count[7]) );
  drp_1 \cache_miss_count_reg[11]  ( .ip(n5200), .ck(clk), .rb(n7950), .q(
        cache_miss_count[11]) );
  drp_1 \cache_hit_count_reg[9]  ( .ip(n5165), .ck(clk), .rb(n7950), .q(
        cache_hit_count[9]) );
  drp_1 \cache_hit_count_reg[8]  ( .ip(n5164), .ck(clk), .rb(n7946), .q(
        cache_hit_count[8]) );
  drp_1 \mem_data_cnt_reg[2]  ( .ip(n7385), .ck(clk), .rb(n7949), .q(
        mem_data_cnt[2]) );
  drp_1 \cache_miss_count_reg[8]  ( .ip(n5197), .ck(clk), .rb(n7948), .q(
        cache_miss_count[8]) );
  drp_1 wr_mem_reg ( .ip(n5256), .ck(clk), .rb(n7949), .q(wr_mem) );
  drp_1 \addr_mem_reg[6]  ( .ip(n5248), .ck(clk), .rb(n7943), .q(addr_mem[6])
         );
  drp_1 \addr_mem_reg[5]  ( .ip(n5249), .ck(clk), .rb(n7949), .q(addr_mem[5])
         );
  drp_1 \addr_mem_reg[4]  ( .ip(n5250), .ck(clk), .rb(n7949), .q(addr_mem[4])
         );
  drp_1 \addr_mem_reg[3]  ( .ip(n5251), .ck(clk), .rb(n7948), .q(addr_mem[3])
         );
  drp_1 \addr_mem_reg[2]  ( .ip(n5252), .ck(clk), .rb(n7943), .q(addr_mem[2])
         );
  drp_1 rd_mem_reg ( .ip(n5255), .ck(clk), .rb(n7949), .q(rd_mem) );
  drp_1 \cache_miss_count_reg[9]  ( .ip(n5198), .ck(clk), .rb(n7943), .q(
        cache_miss_count[9]) );
  drp_1 \mem_data_cnt_reg[3]  ( .ip(n7386), .ck(clk), .rb(n7946), .q(
        mem_data_cnt[3]) );
  drp_1 \cache_miss_count_reg[10]  ( .ip(n5199), .ck(clk), .rb(n7943), .q(
        cache_miss_count[10]) );
  drp_1 \cache_miss_count_reg[13]  ( .ip(n5202), .ck(clk), .rb(n7943), .q(
        cache_miss_count[13]) );
  drp_1 \cache_miss_count_reg[12]  ( .ip(n5201), .ck(clk), .rb(n7944), .q(
        cache_miss_count[12]) );
  drp_1 \cache_hit_count_reg[11]  ( .ip(n5167), .ck(clk), .rb(n7949), .q(
        cache_hit_count[11]) );
  drp_1 \cache_hit_count_reg[10]  ( .ip(n5166), .ck(clk), .rb(n7943), .q(
        cache_hit_count[10]) );
  drp_1 \cache_miss_count_reg[15]  ( .ip(n5204), .ck(clk), .rb(n7946), .q(
        cache_miss_count[15]) );
  drp_1 \cache_miss_count_reg[14]  ( .ip(n5203), .ck(clk), .rb(n7948), .q(
        cache_miss_count[14]) );
  drp_1 \cache_hit_count_reg[13]  ( .ip(n5169), .ck(clk), .rb(n7946), .q(
        cache_hit_count[13]) );
  drp_1 \cache_hit_count_reg[12]  ( .ip(n5168), .ck(clk), .rb(n7946), .q(
        cache_hit_count[12]) );
  drp_1 \cache_miss_count_reg[17]  ( .ip(n5206), .ck(clk), .rb(n7943), .q(
        cache_miss_count[17]) );
  drp_1 \cache_miss_count_reg[16]  ( .ip(n5205), .ck(clk), .rb(n7946), .q(
        cache_miss_count[16]) );
  drp_1 \cache_hit_count_reg[15]  ( .ip(n5171), .ck(clk), .rb(n7946), .q(
        cache_hit_count[15]) );
  drp_1 \cache_hit_count_reg[14]  ( .ip(n5170), .ck(clk), .rb(n7945), .q(
        cache_hit_count[14]) );
  drp_1 \cache_valid_B_reg[3]  ( .ip(n7913), .ck(clk), .rb(n13293), .q(
        cache_valid_B[3]) );
  drp_1 \cache_valid_B_reg[2]  ( .ip(n7914), .ck(clk), .rb(n13293), .q(
        cache_valid_B[2]) );
  drp_1 \cache_valid_B_reg[0]  ( .ip(n7916), .ck(clk), .rb(n13293), .q(
        cache_valid_B[0]) );
  drp_1 \cache_valid_B_reg[4]  ( .ip(n7912), .ck(clk), .rb(n13293), .q(
        cache_valid_B[4]) );
  drp_1 \cache_valid_B_reg[1]  ( .ip(n7915), .ck(clk), .rb(n13293), .q(
        cache_valid_B[1]) );
  drp_1 \cache_valid_B_reg[5]  ( .ip(n7911), .ck(clk), .rb(n13293), .q(
        cache_valid_B[5]) );
  drp_1 \cache_valid_B_reg[6]  ( .ip(n7910), .ck(clk), .rb(n13293), .q(
        cache_valid_B[6]) );
  drp_1 \cache_miss_count_reg[19]  ( .ip(n5208), .ck(clk), .rb(n7948), .q(
        cache_miss_count[19]) );
  drp_1 \cache_valid_A_reg[6]  ( .ip(n7902), .ck(clk), .rb(n7949), .q(
        cache_valid_A[6]) );
  drp_1 \cache_valid_A_reg[0]  ( .ip(n7908), .ck(clk), .rb(n13293), .q(
        cache_valid_A[0]) );
  drp_1 \cache_valid_A_reg[2]  ( .ip(n7906), .ck(clk), .rb(n13293), .q(
        cache_valid_A[2]) );
  drp_1 \cache_valid_A_reg[4]  ( .ip(n7904), .ck(clk), .rb(n7948), .q(
        cache_valid_A[4]) );
  drp_1 \cache_valid_A_reg[1]  ( .ip(n7907), .ck(clk), .rb(n13293), .q(
        cache_valid_A[1]) );
  drp_1 \cache_miss_count_reg[18]  ( .ip(n5207), .ck(clk), .rb(n7947), .q(
        cache_miss_count[18]) );
  drp_1 \cache_valid_A_reg[3]  ( .ip(n7905), .ck(clk), .rb(n13293), .q(
        cache_valid_A[3]) );
  drp_1 \cache_valid_A_reg[5]  ( .ip(n7903), .ck(clk), .rb(n7948), .q(
        cache_valid_A[5]) );
  drp_1 \cache_valid_B_reg[7]  ( .ip(n7909), .ck(clk), .rb(n13293), .q(
        cache_valid_B[7]) );
  drp_1 \cache_hit_count_reg[17]  ( .ip(n5173), .ck(clk), .rb(n7948), .q(
        cache_hit_count[17]) );
  drp_1 \cache_hit_count_reg[16]  ( .ip(n5172), .ck(clk), .rb(n7947), .q(
        cache_hit_count[16]) );
  drp_1 \cache_miss_count_reg[21]  ( .ip(n5210), .ck(clk), .rb(n7944), .q(
        cache_miss_count[21]) );
  drp_1 \cache_miss_count_reg[20]  ( .ip(n5209), .ck(clk), .rb(n7948), .q(
        cache_miss_count[20]) );
  drp_1 \cache_valid_A_reg[7]  ( .ip(n7901), .ck(clk), .rb(n7944), .q(
        cache_valid_A[7]) );
  drp_1 \addr_mem_reg[23]  ( .ip(n5231), .ck(clk), .rb(n7945), .q(addr_mem[23]) );
  drp_1 \addr_mem_reg[29]  ( .ip(n5225), .ck(clk), .rb(n7944), .q(addr_mem[29]) );
  drp_1 \addr_mem_reg[31]  ( .ip(n5223), .ck(clk), .rb(n7944), .q(addr_mem[31]) );
  drp_1 \addr_mem_reg[25]  ( .ip(n5229), .ck(clk), .rb(n7950), .q(addr_mem[25]) );
  drp_1 \addr_mem_reg[30]  ( .ip(n5224), .ck(clk), .rb(n7945), .q(addr_mem[30]) );
  drp_1 \cache_hit_count_reg[19]  ( .ip(n5175), .ck(clk), .rb(n7944), .q(
        cache_hit_count[19]) );
  drp_1 \addr_mem_reg[22]  ( .ip(n5232), .ck(clk), .rb(n7950), .q(addr_mem[22]) );
  drp_1 \addr_mem_reg[13]  ( .ip(n5241), .ck(clk), .rb(n7947), .q(addr_mem[13]) );
  drp_1 \addr_mem_reg[11]  ( .ip(n5243), .ck(clk), .rb(n7945), .q(addr_mem[11]) );
  drp_1 \cache_hit_count_reg[18]  ( .ip(n5174), .ck(clk), .rb(n7945), .q(
        cache_hit_count[18]) );
  drp_1 \addr_mem_reg[7]  ( .ip(n5247), .ck(clk), .rb(n7944), .q(addr_mem[7])
         );
  drp_1 \addr_mem_reg[9]  ( .ip(n5245), .ck(clk), .rb(n7945), .q(addr_mem[9])
         );
  drp_1 \addr_mem_reg[8]  ( .ip(n5246), .ck(clk), .rb(n7945), .q(addr_mem[8])
         );
  drp_1 \addr_mem_reg[28]  ( .ip(n5226), .ck(clk), .rb(n7949), .q(addr_mem[28]) );
  drp_1 \addr_mem_reg[10]  ( .ip(n5244), .ck(clk), .rb(n7947), .q(addr_mem[10]) );
  drp_1 \addr_mem_reg[21]  ( .ip(n5233), .ck(clk), .rb(n7945), .q(addr_mem[21]) );
  drp_1 \addr_mem_reg[12]  ( .ip(n5242), .ck(clk), .rb(n7947), .q(addr_mem[12]) );
  drp_1 \cache_miss_count_reg[23]  ( .ip(n5212), .ck(clk), .rb(n7948), .q(
        cache_miss_count[23]) );
  drp_1 \cache_miss_count_reg[22]  ( .ip(n5211), .ck(clk), .rb(n7947), .q(
        cache_miss_count[22]) );
  drp_1 \addr_mem_reg[19]  ( .ip(n5235), .ck(clk), .rb(n7947), .q(addr_mem[19]) );
  drp_1 \addr_mem_reg[24]  ( .ip(n5230), .ck(clk), .rb(n7943), .q(addr_mem[24]) );
  drp_1 \cache_hit_count_reg[21]  ( .ip(n5177), .ck(clk), .rb(n7950), .q(
        cache_hit_count[21]) );
  drp_1 \cache_hit_count_reg[20]  ( .ip(n5176), .ck(clk), .rb(n7947), .q(
        cache_hit_count[20]) );
  drp_1 \addr_mem_reg[16]  ( .ip(n5238), .ck(clk), .rb(n7950), .q(addr_mem[16]) );
  drp_1 \cache_miss_count_reg[25]  ( .ip(n5214), .ck(clk), .rb(n7949), .q(
        cache_miss_count[25]) );
  drp_1 \cache_miss_count_reg[24]  ( .ip(n5213), .ck(clk), .rb(n7950), .q(
        cache_miss_count[24]) );
  drp_1 \cache_hit_count_reg[23]  ( .ip(n5179), .ck(clk), .rb(n7950), .q(
        cache_hit_count[23]) );
  drp_1 \cache_hit_count_reg[22]  ( .ip(n5178), .ck(clk), .rb(n7946), .q(
        cache_hit_count[22]) );
  drp_1 \cache_miss_count_reg[27]  ( .ip(n5216), .ck(clk), .rb(n7946), .q(
        cache_miss_count[27]) );
  drp_1 \cache_miss_count_reg[26]  ( .ip(n5215), .ck(clk), .rb(n7949), .q(
        cache_miss_count[26]) );
  drp_1 \cache_hit_count_reg[25]  ( .ip(n5181), .ck(clk), .rb(n7944), .q(
        cache_hit_count[25]) );
  drp_1 \cache_hit_count_reg[24]  ( .ip(n5180), .ck(clk), .rb(n7943), .q(
        cache_hit_count[24]) );
  drp_1 \addr_mem_reg[18]  ( .ip(n5236), .ck(clk), .rb(n7949), .q(addr_mem[18]) );
  drp_1 \addr_mem_reg[15]  ( .ip(n5239), .ck(clk), .rb(n7948), .q(addr_mem[15]) );
  drp_1 \addr_mem_reg[14]  ( .ip(n5240), .ck(clk), .rb(n7950), .q(addr_mem[14]) );
  drp_1 \addr_mem_reg[26]  ( .ip(n5228), .ck(clk), .rb(n7949), .q(addr_mem[26]) );
  drp_1 \addr_mem_reg[27]  ( .ip(n5227), .ck(clk), .rb(n7949), .q(addr_mem[27]) );
  drp_1 \cache_miss_count_reg[29]  ( .ip(n5218), .ck(clk), .rb(n7949), .q(
        cache_miss_count[29]) );
  drp_1 \cache_miss_count_reg[28]  ( .ip(n5217), .ck(clk), .rb(n7943), .q(
        cache_miss_count[28]) );
  drp_1 \addr_mem_reg[17]  ( .ip(n5237), .ck(clk), .rb(n7946), .q(addr_mem[17]) );
  drp_1 \addr_mem_reg[20]  ( .ip(n5234), .ck(clk), .rb(n7943), .q(addr_mem[20]) );
  drp_1 \cache_hit_count_reg[27]  ( .ip(n5183), .ck(clk), .rb(n7946), .q(
        cache_hit_count[27]) );
  drp_1 \cache_hit_count_reg[26]  ( .ip(n5182), .ck(clk), .rb(n7943), .q(
        cache_hit_count[26]) );
  drp_1 \cache_miss_count_reg[30]  ( .ip(n5219), .ck(clk), .rb(n7943), .q(
        cache_miss_count[30]) );
  drp_1 \cache_dirty_B_reg[7]  ( .ip(n5329), .ck(clk), .rb(n7944), .q(
        cache_dirty_B[7]) );
  drp_1 \cache_dirty_B_reg[6]  ( .ip(n5330), .ck(clk), .rb(n7946), .q(
        cache_dirty_B[6]) );
  drp_1 \cache_dirty_B_reg[1]  ( .ip(n5335), .ck(clk), .rb(n7943), .q(
        cache_dirty_B[1]) );
  drp_1 \cache_dirty_B_reg[5]  ( .ip(n5331), .ck(clk), .rb(n7946), .q(
        cache_dirty_B[5]) );
  drp_1 \cache_dirty_B_reg[2]  ( .ip(n5334), .ck(clk), .rb(n7948), .q(
        cache_dirty_B[2]) );
  drp_1 \cache_dirty_B_reg[3]  ( .ip(n5333), .ck(clk), .rb(n7946), .q(
        cache_dirty_B[3]) );
  drp_1 \cache_dirty_B_reg[4]  ( .ip(n5332), .ck(clk), .rb(n7946), .q(
        cache_dirty_B[4]) );
  drp_1 \cache_dirty_B_reg[0]  ( .ip(n5336), .ck(clk), .rb(n7945), .q(
        cache_dirty_B[0]) );
  drp_1 \cache_hit_count_reg[29]  ( .ip(n5185), .ck(clk), .rb(n7950), .q(
        cache_hit_count[29]) );
  drp_1 \cache_miss_count_reg[31]  ( .ip(n5220), .ck(clk), .rb(n7948), .q(
        cache_miss_count[31]) );
  drp_1 \cache_hit_count_reg[28]  ( .ip(n5184), .ck(clk), .rb(n7943), .q(
        cache_hit_count[28]) );
  drp_1 hit_reg ( .ip(n5188), .ck(clk), .rb(n7944), .q(hit) );
  drp_1 miss_reg ( .ip(n5221), .ck(clk), .rb(n7948), .q(miss) );
  drp_1 dirty_reg ( .ip(n7941), .ck(clk), .rb(n7947), .q(dirty) );
  drp_1 valid_reg ( .ip(n5155), .ck(clk), .rb(n7946), .q(valid) );
  drp_1 \cache_hit_count_reg[30]  ( .ip(n5186), .ck(clk), .rb(n7948), .q(
        cache_hit_count[30]) );
  drp_1 \cache_dirty_A_reg[0]  ( .ip(n5328), .ck(clk), .rb(n7948), .q(
        cache_dirty_A[0]) );
  drp_1 \cache_dirty_A_reg[7]  ( .ip(n5321), .ck(clk), .rb(n7945), .q(
        cache_dirty_A[7]) );
  drp_1 \cache_dirty_A_reg[6]  ( .ip(n5322), .ck(clk), .rb(n7944), .q(
        cache_dirty_A[6]) );
  drp_1 \cache_dirty_A_reg[2]  ( .ip(n5326), .ck(clk), .rb(n7950), .q(
        cache_dirty_A[2]) );
  drp_1 \cache_dirty_A_reg[1]  ( .ip(n5327), .ck(clk), .rb(n7944), .q(
        cache_dirty_A[1]) );
  drp_1 \cache_dirty_A_reg[5]  ( .ip(n5323), .ck(clk), .rb(n7945), .q(
        cache_dirty_A[5]) );
  drp_1 \cache_dirty_A_reg[4]  ( .ip(n5324), .ck(clk), .rb(n7944), .q(
        cache_dirty_A[4]) );
  drp_1 \cache_dirty_A_reg[3]  ( .ip(n5325), .ck(clk), .rb(n7944), .q(
        cache_dirty_A[3]) );
  drp_1 \cache_hit_count_reg[31]  ( .ip(n5187), .ck(clk), .rb(n7950), .q(
        cache_hit_count[31]) );
  inv_1 U7888 ( .ip(n13297), .op(n7943) );
  inv_1 U7889 ( .ip(n13297), .op(n7944) );
  inv_1 U7890 ( .ip(n13297), .op(n7945) );
  inv_1 U7891 ( .ip(n13297), .op(n7946) );
  inv_1 U7892 ( .ip(n13297), .op(n7947) );
  inv_1 U7893 ( .ip(n13296), .op(n7948) );
  inv_1 U7894 ( .ip(n13297), .op(n7949) );
  inv_1 U7895 ( .ip(n13297), .op(n7950) );
  inv_1 U7897 ( .ip(state[3]), .op(n7956) );
  inv_1 U7898 ( .ip(state[2]), .op(n7962) );
  inv_1 U7899 ( .ip(state[0]), .op(n7989) );
  nand2_1 U7900 ( .ip1(n7962), .ip2(n7989), .op(n7951) );
  nor4_1 U7901 ( .ip1(state[1]), .ip2(state[4]), .ip3(n7956), .ip4(n7951), 
        .op(n7958) );
  nand2_1 U7902 ( .ip1(mem_done), .ip2(n7958), .op(n7954) );
  inv_1 U7903 ( .ip(state[1]), .op(n7952) );
  nor4_1 U7904 ( .ip1(state[3]), .ip2(state[4]), .ip3(n7952), .ip4(n7951), 
        .op(n8620) );
  nand3_1 U7905 ( .ip1(miss), .ip2(valid), .ip3(dirty), .op(n7955) );
  nand4_1 U7906 ( .ip1(hit), .ip2(n8620), .ip3(valid), .ip4(n7955), .op(n7953)
         );
  nand2_1 U7907 ( .ip1(n7954), .ip2(n7953), .op(n13294) );
  inv_1 U7908 ( .ip(busy_mem), .op(n7999) );
  inv_1 U7909 ( .ip(n8620), .op(n9324) );
  nor2_1 U7910 ( .ip1(n9324), .ip2(n7955), .op(n7964) );
  nor2_1 U7911 ( .ip1(state[4]), .ip2(state[1]), .op(n7957) );
  nand2_1 U7912 ( .ip1(n7957), .ip2(n7956), .op(n7988) );
  nor3_1 U7913 ( .ip1(state[0]), .ip2(n7962), .ip3(n7988), .op(n7996) );
  nor2_1 U7914 ( .ip1(n7958), .ip2(n7996), .op(n9323) );
  nor2_1 U7915 ( .ip1(mem_done), .ip2(n9323), .op(n7961) );
  nand2_1 U7916 ( .ip1(n8620), .ip2(valid), .op(n7959) );
  nor3_1 U7917 ( .ip1(miss), .ip2(n7959), .ip3(hit), .op(n7960) );
  nor2_1 U7918 ( .ip1(n7961), .ip2(n7960), .op(n7991) );
  nor2_1 U7919 ( .ip1(n7991), .ip2(n7962), .op(n7963) );
  or2_1 U7920 ( .ip1(n7964), .ip2(n7963), .op(next_state[2]) );
  nand2_1 U7921 ( .ip1(n7999), .ip2(next_state[2]), .op(n13189) );
  nor2_1 U7922 ( .ip1(SelectWay), .ip2(n13189), .op(n8555) );
  nor2_1 U7923 ( .ip1(addr_resp[6]), .ip2(addr_resp[5]), .op(n7965) );
  inv_1 U7924 ( .ip(addr_resp[4]), .op(n7974) );
  nand2_1 U7925 ( .ip1(n7965), .ip2(n7974), .op(n9860) );
  inv_1 U7926 ( .ip(n9860), .op(n12370) );
  buf_1 U7927 ( .ip(n12370), .op(n12204) );
  nand2_1 U7928 ( .ip1(\cache_tag_A[0][14] ), .ip2(n12204), .op(n7977) );
  inv_1 U7929 ( .ip(addr_resp[6]), .op(n7973) );
  inv_1 U7930 ( .ip(addr_resp[5]), .op(n7966) );
  nor3_1 U7931 ( .ip1(n7974), .ip2(n7973), .ip3(n7966), .op(n12278) );
  nand3_1 U7932 ( .ip1(n7973), .ip2(addr_resp[4]), .ip3(addr_resp[5]), .op(
        n9866) );
  inv_1 U7933 ( .ip(\cache_tag_A[3][14] ), .op(n8938) );
  nor2_1 U7934 ( .ip1(n9866), .ip2(n8938), .op(n7972) );
  nand3_1 U7935 ( .ip1(n7974), .ip2(n7966), .ip3(addr_resp[6]), .op(n9868) );
  inv_1 U7936 ( .ip(n9868), .op(n12054) );
  buf_1 U7937 ( .ip(n12054), .op(n12396) );
  nand2_1 U7938 ( .ip1(n11156), .ip2(\cache_tag_A[4][14] ), .op(n7970) );
  nand3_1 U7939 ( .ip1(n7966), .ip2(addr_resp[6]), .ip3(addr_resp[4]), .op(
        n9870) );
  inv_1 U7940 ( .ip(n9870), .op(n11236) );
  buf_1 U7941 ( .ip(n11236), .op(n12582) );
  buf_1 U7942 ( .ip(n12582), .op(n12256) );
  buf_1 U7943 ( .ip(n12256), .op(n12118) );
  nand2_1 U7944 ( .ip1(n12118), .ip2(\cache_tag_A[5][14] ), .op(n7969) );
  nand3_1 U7945 ( .ip1(n7973), .ip2(n7966), .ip3(addr_resp[4]), .op(n9862) );
  inv_1 U7946 ( .ip(n9862), .op(n11724) );
  buf_1 U7947 ( .ip(n11724), .op(n12147) );
  nand2_1 U7948 ( .ip1(n12147), .ip2(\cache_tag_A[1][14] ), .op(n7968) );
  nor3_1 U7949 ( .ip1(n7973), .ip2(n7966), .ip3(addr_resp[4]), .op(n12429) );
  buf_1 U7950 ( .ip(n12429), .op(n11780) );
  nand2_1 U7951 ( .ip1(n11780), .ip2(\cache_tag_A[6][14] ), .op(n7967) );
  nand4_1 U7952 ( .ip1(n7970), .ip2(n7969), .ip3(n7968), .ip4(n7967), .op(
        n7971) );
  not_ab_or_c_or_d U7953 ( .ip1(\cache_tag_A[7][14] ), .ip2(n11057), .ip3(
        n7972), .ip4(n7971), .op(n7976) );
  nand3_1 U7954 ( .ip1(n7974), .ip2(n7973), .ip3(addr_resp[5]), .op(n9864) );
  inv_1 U7955 ( .ip(n9864), .op(n12546) );
  buf_1 U7956 ( .ip(n12546), .op(n11855) );
  nand2_1 U7957 ( .ip1(n11855), .ip2(\cache_tag_A[2][14] ), .op(n7975) );
  nand3_1 U7958 ( .ip1(n7977), .ip2(n7976), .ip3(n7975), .op(n9464) );
  nand2_1 U7959 ( .ip1(n8555), .ip2(n9464), .op(n8003) );
  inv_1 U7960 ( .ip(SelectWay), .op(n9702) );
  nor2_1 U7961 ( .ip1(n9702), .ip2(n13189), .op(n8545) );
  buf_1 U7962 ( .ip(n12546), .op(n12583) );
  nand2_1 U7963 ( .ip1(n12583), .ip2(\cache_tag_B[2][14] ), .op(n7986) );
  buf_1 U7964 ( .ip(n11724), .op(n11946) );
  inv_1 U7965 ( .ip(\cache_tag_B[5][14] ), .op(n9163) );
  nor2_1 U7966 ( .ip1(n9870), .ip2(n9163), .op(n7983) );
  nand2_1 U7967 ( .ip1(n12396), .ip2(\cache_tag_B[4][14] ), .op(n7981) );
  inv_1 U7968 ( .ip(n9866), .op(n12559) );
  buf_1 U7969 ( .ip(n12559), .op(n12410) );
  buf_1 U7970 ( .ip(n12410), .op(n12591) );
  nand2_1 U7971 ( .ip1(n12591), .ip2(\cache_tag_B[3][14] ), .op(n7980) );
  buf_1 U7972 ( .ip(n12429), .op(n12551) );
  nand2_1 U7973 ( .ip1(n12551), .ip2(\cache_tag_B[6][14] ), .op(n7979) );
  nand2_1 U7974 ( .ip1(n12370), .ip2(\cache_tag_B[0][14] ), .op(n7978) );
  nand4_1 U7975 ( .ip1(n7981), .ip2(n7980), .ip3(n7979), .ip4(n7978), .op(
        n7982) );
  not_ab_or_c_or_d U7976 ( .ip1(\cache_tag_B[1][14] ), .ip2(n11946), .ip3(
        n7983), .ip4(n7982), .op(n7985) );
  nand2_1 U7977 ( .ip1(n10575), .ip2(\cache_tag_B[7][14] ), .op(n7984) );
  nand3_1 U7978 ( .ip1(n7986), .ip2(n7985), .ip3(n7984), .op(n7987) );
  nand2_1 U7979 ( .ip1(n8545), .ip2(n7987), .op(n8002) );
  inv_1 U7980 ( .ip(n13294), .op(n9544) );
  nor2_1 U7981 ( .ip1(wr), .ip2(rd), .op(n9363) );
  nor3_1 U7982 ( .ip1(state[2]), .ip2(n7989), .ip3(n7988), .op(n7990) );
  inv_1 U7983 ( .ip(n7990), .op(n9322) );
  nor2_1 U7984 ( .ip1(n9363), .ip2(n9322), .op(n9320) );
  inv_1 U7985 ( .ip(n9320), .op(n13290) );
  nand2_1 U7986 ( .ip1(n9363), .ip2(n7990), .op(n9325) );
  nand2_1 U7987 ( .ip1(n7991), .ip2(n9325), .op(n7995) );
  nand2_1 U7988 ( .ip1(state[1]), .ip2(n7995), .op(n7992) );
  nand2_1 U7989 ( .ip1(n13290), .ip2(n7992), .op(next_state[1]) );
  inv_1 U7990 ( .ip(next_state[1]), .op(n9362) );
  nand2_1 U7991 ( .ip1(n9544), .ip2(n9362), .op(n13201) );
  nand2_1 U7992 ( .ip1(addr_mem[21]), .ip2(n13201), .op(n8001) );
  nand2_1 U7993 ( .ip1(n8620), .ip2(miss), .op(n13231) );
  nor3_1 U7994 ( .ip1(hit), .ip2(dirty), .ip3(n13231), .op(n7994) );
  nor2_1 U7995 ( .ip1(valid), .ip2(n9324), .op(n7993) );
  not_ab_or_c_or_d U7996 ( .ip1(state[3]), .ip2(n7995), .ip3(n7994), .ip4(
        n7993), .op(n7998) );
  nand2_1 U7997 ( .ip1(mem_done), .ip2(n7996), .op(n7997) );
  nand2_1 U7998 ( .ip1(n7998), .ip2(n7997), .op(n13295) );
  nand2_1 U7999 ( .ip1(n13295), .ip2(n7999), .op(n13191) );
  inv_1 U8000 ( .ip(n13191), .op(n9703) );
  nand2_1 U8001 ( .ip1(addr_resp[21]), .ip2(n9703), .op(n8000) );
  nand4_1 U8002 ( .ip1(n8003), .ip2(n8002), .ip3(n8001), .ip4(n8000), .op(
        n5233) );
  nand2_1 U8003 ( .ip1(addr_mem[9]), .ip2(n13201), .op(n8026) );
  buf_1 U8004 ( .ip(n12429), .op(n12458) );
  nand2_1 U8005 ( .ip1(n12458), .ip2(\cache_tag_A[6][2] ), .op(n8012) );
  inv_1 U8006 ( .ip(\cache_tag_A[5][2] ), .op(n8960) );
  nor2_1 U8007 ( .ip1(n9870), .ip2(n8960), .op(n8009) );
  buf_1 U8008 ( .ip(n12546), .op(n10426) );
  nand2_1 U8009 ( .ip1(n10426), .ip2(\cache_tag_A[2][2] ), .op(n8007) );
  nand2_1 U8010 ( .ip1(n12370), .ip2(\cache_tag_A[0][2] ), .op(n8006) );
  buf_1 U8011 ( .ip(n12559), .op(n8060) );
  buf_1 U8012 ( .ip(n8060), .op(n11535) );
  nand2_1 U8013 ( .ip1(n11535), .ip2(\cache_tag_A[3][2] ), .op(n8005) );
  buf_1 U8014 ( .ip(n11724), .op(n10166) );
  nand2_1 U8015 ( .ip1(n10166), .ip2(\cache_tag_A[1][2] ), .op(n8004) );
  nand4_1 U8016 ( .ip1(n8007), .ip2(n8006), .ip3(n8005), .ip4(n8004), .op(
        n8008) );
  not_ab_or_c_or_d U8017 ( .ip1(\cache_tag_A[7][2] ), .ip2(n10702), .ip3(n8009), .ip4(n8008), .op(n8011) );
  buf_1 U8018 ( .ip(n12054), .op(n11156) );
  buf_1 U8019 ( .ip(n11156), .op(n11324) );
  nand2_1 U8020 ( .ip1(n11324), .ip2(\cache_tag_A[4][2] ), .op(n8010) );
  nand3_1 U8021 ( .ip1(n8012), .ip2(n8011), .ip3(n8010), .op(n9526) );
  nand2_1 U8022 ( .ip1(n8555), .ip2(n9526), .op(n8025) );
  nand2_1 U8023 ( .ip1(n12357), .ip2(\cache_tag_B[0][2] ), .op(n8021) );
  inv_1 U8024 ( .ip(\cache_tag_B[3][2] ), .op(n9218) );
  nor2_1 U8025 ( .ip1(n9866), .ip2(n9218), .op(n8018) );
  nand2_1 U8026 ( .ip1(n12551), .ip2(\cache_tag_B[6][2] ), .op(n8016) );
  buf_1 U8027 ( .ip(n11156), .op(n12584) );
  nand2_1 U8028 ( .ip1(n12584), .ip2(\cache_tag_B[4][2] ), .op(n8015) );
  nand2_1 U8029 ( .ip1(n10686), .ip2(\cache_tag_B[1][2] ), .op(n8014) );
  nand2_1 U8030 ( .ip1(n12583), .ip2(\cache_tag_B[2][2] ), .op(n8013) );
  nand4_1 U8031 ( .ip1(n8016), .ip2(n8015), .ip3(n8014), .ip4(n8013), .op(
        n8017) );
  not_ab_or_c_or_d U8032 ( .ip1(\cache_tag_B[5][2] ), .ip2(n11236), .ip3(n8018), .ip4(n8017), .op(n8020) );
  nand2_1 U8033 ( .ip1(n11057), .ip2(\cache_tag_B[7][2] ), .op(n8019) );
  nand3_1 U8034 ( .ip1(n8021), .ip2(n8020), .ip3(n8019), .op(n8022) );
  nand2_1 U8035 ( .ip1(n8545), .ip2(n8022), .op(n8024) );
  nand2_1 U8036 ( .ip1(addr_resp[9]), .ip2(n9703), .op(n8023) );
  nand4_1 U8037 ( .ip1(n8026), .ip2(n8025), .ip3(n8024), .ip4(n8023), .op(
        n5245) );
  nand2_1 U8038 ( .ip1(n12370), .ip2(\cache_tag_B[0][6] ), .op(n8035) );
  inv_1 U8039 ( .ip(n12278), .op(n9769) );
  inv_1 U8040 ( .ip(\cache_tag_B[7][6] ), .op(n9043) );
  nor2_1 U8041 ( .ip1(n9769), .ip2(n9043), .op(n8032) );
  nand2_1 U8042 ( .ip1(n12583), .ip2(\cache_tag_B[2][6] ), .op(n8030) );
  nand2_1 U8043 ( .ip1(n12584), .ip2(\cache_tag_B[4][6] ), .op(n8029) );
  nand2_1 U8044 ( .ip1(n12118), .ip2(\cache_tag_B[5][6] ), .op(n8028) );
  nand2_1 U8045 ( .ip1(n12551), .ip2(\cache_tag_B[6][6] ), .op(n8027) );
  nand4_1 U8046 ( .ip1(n8030), .ip2(n8029), .ip3(n8028), .ip4(n8027), .op(
        n8031) );
  not_ab_or_c_or_d U8047 ( .ip1(\cache_tag_B[3][6] ), .ip2(n8060), .ip3(n8032), 
        .ip4(n8031), .op(n8034) );
  nand2_1 U8048 ( .ip1(n10686), .ip2(\cache_tag_B[1][6] ), .op(n8033) );
  nand3_1 U8049 ( .ip1(n8035), .ip2(n8034), .ip3(n8033), .op(n8036) );
  nand2_1 U8050 ( .ip1(n8545), .ip2(n8036), .op(n8049) );
  buf_1 U8051 ( .ip(n12396), .op(n12476) );
  buf_1 U8052 ( .ip(n12476), .op(n12194) );
  nand2_1 U8053 ( .ip1(\cache_tag_A[4][6] ), .ip2(n12194), .op(n8045) );
  buf_1 U8054 ( .ip(n12370), .op(n12297) );
  inv_1 U8055 ( .ip(\cache_tag_A[1][6] ), .op(n8703) );
  nor2_1 U8056 ( .ip1(n9862), .ip2(n8703), .op(n8042) );
  nand2_1 U8057 ( .ip1(n11535), .ip2(\cache_tag_A[3][6] ), .op(n8040) );
  nand2_1 U8058 ( .ip1(n12458), .ip2(\cache_tag_A[6][6] ), .op(n8039) );
  buf_1 U8059 ( .ip(n12278), .op(n10575) );
  nand2_1 U8060 ( .ip1(n10575), .ip2(\cache_tag_A[7][6] ), .op(n8038) );
  nand2_1 U8061 ( .ip1(n10426), .ip2(\cache_tag_A[2][6] ), .op(n8037) );
  nand4_1 U8062 ( .ip1(n8040), .ip2(n8039), .ip3(n8038), .ip4(n8037), .op(
        n8041) );
  not_ab_or_c_or_d U8063 ( .ip1(n12297), .ip2(\cache_tag_A[0][6] ), .ip3(n8042), .ip4(n8041), .op(n8044) );
  buf_1 U8064 ( .ip(n11236), .op(n11296) );
  buf_1 U8065 ( .ip(n11296), .op(n11304) );
  nand2_1 U8066 ( .ip1(n11304), .ip2(\cache_tag_A[5][6] ), .op(n8043) );
  nand3_1 U8067 ( .ip1(n8045), .ip2(n8044), .ip3(n8043), .op(n9528) );
  nand2_1 U8068 ( .ip1(n8555), .ip2(n9528), .op(n8048) );
  nand2_1 U8069 ( .ip1(addr_mem[13]), .ip2(n13201), .op(n8047) );
  buf_1 U8070 ( .ip(n9703), .op(n9619) );
  nand2_1 U8071 ( .ip1(addr_resp[13]), .ip2(n9619), .op(n8046) );
  nand4_1 U8072 ( .ip1(n8049), .ip2(n8048), .ip3(n8047), .ip4(n8046), .op(
        n5241) );
  buf_1 U8073 ( .ip(n12429), .op(n12320) );
  nand2_1 U8074 ( .ip1(n12320), .ip2(\cache_tag_B[6][16] ), .op(n8058) );
  inv_1 U8075 ( .ip(\cache_tag_B[7][16] ), .op(n9103) );
  nor2_1 U8076 ( .ip1(n9769), .ip2(n9103), .op(n8055) );
  buf_1 U8077 ( .ip(n12410), .op(n12321) );
  nand2_1 U8078 ( .ip1(n12321), .ip2(\cache_tag_B[3][16] ), .op(n8053) );
  nand2_1 U8079 ( .ip1(n12256), .ip2(\cache_tag_B[5][16] ), .op(n8052) );
  nand2_1 U8080 ( .ip1(n12370), .ip2(\cache_tag_B[0][16] ), .op(n8051) );
  nand2_1 U8081 ( .ip1(n12583), .ip2(\cache_tag_B[2][16] ), .op(n8050) );
  nand4_1 U8082 ( .ip1(n8053), .ip2(n8052), .ip3(n8051), .ip4(n8050), .op(
        n8054) );
  not_ab_or_c_or_d U8083 ( .ip1(\cache_tag_B[1][16] ), .ip2(n11946), .ip3(
        n8055), .ip4(n8054), .op(n8057) );
  nand2_1 U8084 ( .ip1(n12396), .ip2(\cache_tag_B[4][16] ), .op(n8056) );
  nand3_1 U8085 ( .ip1(n8058), .ip2(n8057), .ip3(n8056), .op(n8059) );
  nand2_1 U8086 ( .ip1(n8545), .ip2(n8059), .op(n8073) );
  buf_1 U8087 ( .ip(n12546), .op(n12486) );
  nand2_1 U8088 ( .ip1(\cache_tag_A[2][16] ), .ip2(n12486), .op(n8069) );
  buf_1 U8089 ( .ip(n8060), .op(n12096) );
  inv_1 U8090 ( .ip(\cache_tag_A[5][16] ), .op(n8874) );
  nor2_1 U8091 ( .ip1(n9870), .ip2(n8874), .op(n8066) );
  buf_1 U8092 ( .ip(n12370), .op(n8452) );
  nand2_1 U8093 ( .ip1(n8452), .ip2(\cache_tag_A[0][16] ), .op(n8064) );
  buf_1 U8094 ( .ip(n12429), .op(n12371) );
  nand2_1 U8095 ( .ip1(n12371), .ip2(\cache_tag_A[6][16] ), .op(n8063) );
  buf_1 U8096 ( .ip(n12278), .op(n11057) );
  nand2_1 U8097 ( .ip1(n11057), .ip2(\cache_tag_A[7][16] ), .op(n8062) );
  nand2_1 U8098 ( .ip1(n10166), .ip2(\cache_tag_A[1][16] ), .op(n8061) );
  nand4_1 U8099 ( .ip1(n8064), .ip2(n8063), .ip3(n8062), .ip4(n8061), .op(
        n8065) );
  not_ab_or_c_or_d U8100 ( .ip1(\cache_tag_A[3][16] ), .ip2(n12096), .ip3(
        n8066), .ip4(n8065), .op(n8068) );
  nand2_1 U8101 ( .ip1(n11324), .ip2(\cache_tag_A[4][16] ), .op(n8067) );
  nand3_1 U8102 ( .ip1(n8069), .ip2(n8068), .ip3(n8067), .op(n9502) );
  nand2_1 U8103 ( .ip1(n8555), .ip2(n9502), .op(n8072) );
  nand2_1 U8104 ( .ip1(addr_mem[23]), .ip2(n13201), .op(n8071) );
  nand2_1 U8105 ( .ip1(addr_resp[23]), .ip2(n9703), .op(n8070) );
  nand4_1 U8106 ( .ip1(n8073), .ip2(n8072), .ip3(n8071), .ip4(n8070), .op(
        n5231) );
  nand2_1 U8107 ( .ip1(addr_mem[31]), .ip2(n13201), .op(n8096) );
  nand2_1 U8108 ( .ip1(n12583), .ip2(\cache_tag_A[2][24] ), .op(n8082) );
  inv_1 U8109 ( .ip(\cache_tag_A[1][24] ), .op(n8900) );
  nor2_1 U8110 ( .ip1(n9862), .ip2(n8900), .op(n8079) );
  nand2_1 U8111 ( .ip1(n11057), .ip2(\cache_tag_A[7][24] ), .op(n8077) );
  nand2_1 U8112 ( .ip1(n12371), .ip2(\cache_tag_A[6][24] ), .op(n8076) );
  nand2_1 U8113 ( .ip1(n11535), .ip2(\cache_tag_A[3][24] ), .op(n8075) );
  nand2_1 U8114 ( .ip1(n8452), .ip2(\cache_tag_A[0][24] ), .op(n8074) );
  nand4_1 U8115 ( .ip1(n8077), .ip2(n8076), .ip3(n8075), .ip4(n8074), .op(
        n8078) );
  not_ab_or_c_or_d U8116 ( .ip1(\cache_tag_A[4][24] ), .ip2(n11156), .ip3(
        n8079), .ip4(n8078), .op(n8081) );
  nand2_1 U8117 ( .ip1(n11304), .ip2(\cache_tag_A[5][24] ), .op(n8080) );
  nand3_1 U8118 ( .ip1(n8082), .ip2(n8081), .ip3(n8080), .op(n9504) );
  nand2_1 U8119 ( .ip1(n8555), .ip2(n9504), .op(n8095) );
  nand2_1 U8120 ( .ip1(n12371), .ip2(\cache_tag_B[6][24] ), .op(n8091) );
  inv_1 U8121 ( .ip(\cache_tag_B[7][24] ), .op(n9140) );
  nor2_1 U8122 ( .ip1(n9769), .ip2(n9140), .op(n8088) );
  nand2_1 U8123 ( .ip1(n12321), .ip2(\cache_tag_B[3][24] ), .op(n8086) );
  nand2_1 U8124 ( .ip1(n12583), .ip2(\cache_tag_B[2][24] ), .op(n8085) );
  nand2_1 U8125 ( .ip1(n12370), .ip2(\cache_tag_B[0][24] ), .op(n8084) );
  nand2_1 U8126 ( .ip1(n11324), .ip2(\cache_tag_B[4][24] ), .op(n8083) );
  nand4_1 U8127 ( .ip1(n8086), .ip2(n8085), .ip3(n8084), .ip4(n8083), .op(
        n8087) );
  not_ab_or_c_or_d U8128 ( .ip1(\cache_tag_B[5][24] ), .ip2(n11296), .ip3(
        n8088), .ip4(n8087), .op(n8090) );
  nand2_1 U8129 ( .ip1(n10166), .ip2(\cache_tag_B[1][24] ), .op(n8089) );
  nand3_1 U8130 ( .ip1(n8091), .ip2(n8090), .ip3(n8089), .op(n8092) );
  nand2_1 U8131 ( .ip1(n8545), .ip2(n8092), .op(n8094) );
  nand2_1 U8132 ( .ip1(addr_resp[31]), .ip2(n9619), .op(n8093) );
  nand4_1 U8133 ( .ip1(n8096), .ip2(n8095), .ip3(n8094), .ip4(n8093), .op(
        n5223) );
  nand2_1 U8134 ( .ip1(n12320), .ip2(\cache_tag_B[6][15] ), .op(n8105) );
  buf_1 U8135 ( .ip(n12546), .op(n12475) );
  inv_1 U8136 ( .ip(\cache_tag_B[7][15] ), .op(n9206) );
  nor2_1 U8137 ( .ip1(n9769), .ip2(n9206), .op(n8102) );
  nand2_1 U8138 ( .ip1(n12370), .ip2(\cache_tag_B[0][15] ), .op(n8100) );
  nand2_1 U8139 ( .ip1(n12591), .ip2(\cache_tag_B[3][15] ), .op(n8099) );
  nand2_1 U8140 ( .ip1(n10686), .ip2(\cache_tag_B[1][15] ), .op(n8098) );
  nand2_1 U8141 ( .ip1(n12256), .ip2(\cache_tag_B[5][15] ), .op(n8097) );
  nand4_1 U8142 ( .ip1(n8100), .ip2(n8099), .ip3(n8098), .ip4(n8097), .op(
        n8101) );
  not_ab_or_c_or_d U8143 ( .ip1(\cache_tag_B[2][15] ), .ip2(n12475), .ip3(
        n8102), .ip4(n8101), .op(n8104) );
  nand2_1 U8144 ( .ip1(n12396), .ip2(\cache_tag_B[4][15] ), .op(n8103) );
  nand3_1 U8145 ( .ip1(n8105), .ip2(n8104), .ip3(n8103), .op(n8106) );
  nand2_1 U8146 ( .ip1(n8545), .ip2(n8106), .op(n8119) );
  buf_1 U8147 ( .ip(n12278), .op(n10702) );
  nand2_1 U8148 ( .ip1(n10702), .ip2(\cache_tag_A[7][15] ), .op(n8115) );
  inv_1 U8149 ( .ip(\cache_tag_A[3][15] ), .op(n8777) );
  nor2_1 U8150 ( .ip1(n9866), .ip2(n8777), .op(n8112) );
  nand2_1 U8151 ( .ip1(n11304), .ip2(\cache_tag_A[5][15] ), .op(n8110) );
  nand2_1 U8152 ( .ip1(n11724), .ip2(\cache_tag_A[1][15] ), .op(n8109) );
  nand2_1 U8153 ( .ip1(n12370), .ip2(\cache_tag_A[0][15] ), .op(n8108) );
  nand2_1 U8154 ( .ip1(n11324), .ip2(\cache_tag_A[4][15] ), .op(n8107) );
  nand4_1 U8155 ( .ip1(n8110), .ip2(n8109), .ip3(n8108), .ip4(n8107), .op(
        n8111) );
  not_ab_or_c_or_d U8156 ( .ip1(\cache_tag_A[2][15] ), .ip2(n12475), .ip3(
        n8112), .ip4(n8111), .op(n8114) );
  nand2_1 U8157 ( .ip1(n12458), .ip2(\cache_tag_A[6][15] ), .op(n8113) );
  nand3_1 U8158 ( .ip1(n8115), .ip2(n8114), .ip3(n8113), .op(n9518) );
  nand2_1 U8159 ( .ip1(n8555), .ip2(n9518), .op(n8118) );
  nand2_1 U8160 ( .ip1(addr_mem[22]), .ip2(n13201), .op(n8117) );
  nand2_1 U8161 ( .ip1(addr_resp[22]), .ip2(n9703), .op(n8116) );
  nand4_1 U8162 ( .ip1(n8119), .ip2(n8118), .ip3(n8117), .ip4(n8116), .op(
        n5232) );
  nand2_1 U8163 ( .ip1(addr_mem[29]), .ip2(n13201), .op(n8142) );
  nand2_1 U8164 ( .ip1(n12370), .ip2(\cache_tag_B[0][22] ), .op(n8128) );
  inv_1 U8165 ( .ip(\cache_tag_B[7][22] ), .op(n9295) );
  nor2_1 U8166 ( .ip1(n9769), .ip2(n9295), .op(n8125) );
  nand2_1 U8167 ( .ip1(n12371), .ip2(\cache_tag_B[6][22] ), .op(n8123) );
  nand2_1 U8168 ( .ip1(n12256), .ip2(\cache_tag_B[5][22] ), .op(n8122) );
  nand2_1 U8169 ( .ip1(n10166), .ip2(\cache_tag_B[1][22] ), .op(n8121) );
  nand2_1 U8170 ( .ip1(n12321), .ip2(\cache_tag_B[3][22] ), .op(n8120) );
  nand4_1 U8171 ( .ip1(n8123), .ip2(n8122), .ip3(n8121), .ip4(n8120), .op(
        n8124) );
  not_ab_or_c_or_d U8172 ( .ip1(\cache_tag_B[2][22] ), .ip2(n12475), .ip3(
        n8125), .ip4(n8124), .op(n8127) );
  nand2_1 U8173 ( .ip1(n11324), .ip2(\cache_tag_B[4][22] ), .op(n8126) );
  nand3_1 U8174 ( .ip1(n8128), .ip2(n8127), .ip3(n8126), .op(n8129) );
  nand2_1 U8175 ( .ip1(n8545), .ip2(n8129), .op(n8141) );
  nand2_1 U8176 ( .ip1(n12458), .ip2(\cache_tag_A[6][22] ), .op(n8138) );
  inv_1 U8177 ( .ip(\cache_tag_A[5][22] ), .op(n8692) );
  nor2_1 U8178 ( .ip1(n9870), .ip2(n8692), .op(n8135) );
  nand2_1 U8179 ( .ip1(n12583), .ip2(\cache_tag_A[2][22] ), .op(n8133) );
  nand2_1 U8180 ( .ip1(n10702), .ip2(\cache_tag_A[7][22] ), .op(n8132) );
  nand2_1 U8181 ( .ip1(n8452), .ip2(\cache_tag_A[0][22] ), .op(n8131) );
  nand2_1 U8182 ( .ip1(n11535), .ip2(\cache_tag_A[3][22] ), .op(n8130) );
  nand4_1 U8183 ( .ip1(n8133), .ip2(n8132), .ip3(n8131), .ip4(n8130), .op(
        n8134) );
  not_ab_or_c_or_d U8184 ( .ip1(n11156), .ip2(\cache_tag_A[4][22] ), .ip3(
        n8135), .ip4(n8134), .op(n8137) );
  nand2_1 U8185 ( .ip1(n10166), .ip2(\cache_tag_A[1][22] ), .op(n8136) );
  nand3_1 U8186 ( .ip1(n8138), .ip2(n8137), .ip3(n8136), .op(n9514) );
  nand2_1 U8187 ( .ip1(n8555), .ip2(n9514), .op(n8140) );
  nand2_1 U8188 ( .ip1(addr_resp[29]), .ip2(n9703), .op(n8139) );
  nand4_1 U8189 ( .ip1(n8142), .ip2(n8141), .ip3(n8140), .ip4(n8139), .op(
        n5225) );
  nand2_1 U8190 ( .ip1(addr_mem[11]), .ip2(n13201), .op(n8165) );
  nand2_1 U8191 ( .ip1(\cache_tag_A[4][4] ), .ip2(n12194), .op(n8151) );
  inv_1 U8192 ( .ip(\cache_tag_A[3][4] ), .op(n8715) );
  nor2_1 U8193 ( .ip1(n9866), .ip2(n8715), .op(n8148) );
  nand2_1 U8194 ( .ip1(n11304), .ip2(\cache_tag_A[5][4] ), .op(n8146) );
  nand2_1 U8195 ( .ip1(n12583), .ip2(\cache_tag_A[2][4] ), .op(n8145) );
  nand2_1 U8196 ( .ip1(n12371), .ip2(\cache_tag_A[6][4] ), .op(n8144) );
  nand2_1 U8197 ( .ip1(n11057), .ip2(\cache_tag_A[7][4] ), .op(n8143) );
  nand4_1 U8198 ( .ip1(n8146), .ip2(n8145), .ip3(n8144), .ip4(n8143), .op(
        n8147) );
  not_ab_or_c_or_d U8199 ( .ip1(n12297), .ip2(\cache_tag_A[0][4] ), .ip3(n8148), .ip4(n8147), .op(n8150) );
  nand2_1 U8200 ( .ip1(n10166), .ip2(\cache_tag_A[1][4] ), .op(n8149) );
  nand3_1 U8201 ( .ip1(n8151), .ip2(n8150), .ip3(n8149), .op(n9506) );
  nand2_1 U8202 ( .ip1(n8555), .ip2(n9506), .op(n8164) );
  nand2_1 U8203 ( .ip1(n12583), .ip2(\cache_tag_B[2][4] ), .op(n8160) );
  buf_1 U8204 ( .ip(n12370), .op(n12357) );
  inv_1 U8205 ( .ip(\cache_tag_B[7][4] ), .op(n9054) );
  nor2_1 U8206 ( .ip1(n9769), .ip2(n9054), .op(n8157) );
  nand2_1 U8207 ( .ip1(n11946), .ip2(\cache_tag_B[1][4] ), .op(n8155) );
  nand2_1 U8208 ( .ip1(n12118), .ip2(\cache_tag_B[5][4] ), .op(n8154) );
  nand2_1 U8209 ( .ip1(n12591), .ip2(\cache_tag_B[3][4] ), .op(n8153) );
  nand2_1 U8210 ( .ip1(n12584), .ip2(\cache_tag_B[4][4] ), .op(n8152) );
  nand4_1 U8211 ( .ip1(n8155), .ip2(n8154), .ip3(n8153), .ip4(n8152), .op(
        n8156) );
  not_ab_or_c_or_d U8212 ( .ip1(\cache_tag_B[0][4] ), .ip2(n12357), .ip3(n8157), .ip4(n8156), .op(n8159) );
  nand2_1 U8213 ( .ip1(n12551), .ip2(\cache_tag_B[6][4] ), .op(n8158) );
  nand3_1 U8214 ( .ip1(n8160), .ip2(n8159), .ip3(n8158), .op(n8161) );
  nand2_1 U8215 ( .ip1(n8545), .ip2(n8161), .op(n8163) );
  nand2_1 U8216 ( .ip1(addr_resp[11]), .ip2(n9703), .op(n8162) );
  nand4_1 U8217 ( .ip1(n8165), .ip2(n8164), .ip3(n8163), .ip4(n8162), .op(
        n5243) );
  nand2_1 U8218 ( .ip1(n12321), .ip2(\cache_tag_A[3][18] ), .op(n8174) );
  inv_1 U8219 ( .ip(\cache_tag_A[4][18] ), .op(n8840) );
  nor2_1 U8220 ( .ip1(n9868), .ip2(n8840), .op(n8171) );
  nand2_1 U8221 ( .ip1(n12371), .ip2(\cache_tag_A[6][18] ), .op(n8169) );
  nand2_1 U8222 ( .ip1(n11057), .ip2(\cache_tag_A[7][18] ), .op(n8168) );
  nand2_1 U8223 ( .ip1(n12583), .ip2(\cache_tag_A[2][18] ), .op(n8167) );
  nand2_1 U8224 ( .ip1(n12256), .ip2(\cache_tag_A[5][18] ), .op(n8166) );
  nand4_1 U8225 ( .ip1(n8169), .ip2(n8168), .ip3(n8167), .ip4(n8166), .op(
        n8170) );
  not_ab_or_c_or_d U8226 ( .ip1(\cache_tag_A[0][18] ), .ip2(n12357), .ip3(
        n8171), .ip4(n8170), .op(n8173) );
  nand2_1 U8227 ( .ip1(n10166), .ip2(\cache_tag_A[1][18] ), .op(n8172) );
  nand3_1 U8228 ( .ip1(n8174), .ip2(n8173), .ip3(n8172), .op(n9474) );
  nand2_1 U8229 ( .ip1(n8555), .ip2(n9474), .op(n8188) );
  nand2_1 U8230 ( .ip1(n12370), .ip2(\cache_tag_B[0][18] ), .op(n8183) );
  inv_1 U8231 ( .ip(\cache_tag_B[7][18] ), .op(n9028) );
  nor2_1 U8232 ( .ip1(n9769), .ip2(n9028), .op(n8180) );
  nand2_1 U8233 ( .ip1(n12583), .ip2(\cache_tag_B[2][18] ), .op(n8178) );
  nand2_1 U8234 ( .ip1(n12551), .ip2(\cache_tag_B[6][18] ), .op(n8177) );
  nand2_1 U8235 ( .ip1(n11946), .ip2(\cache_tag_B[1][18] ), .op(n8176) );
  nand2_1 U8236 ( .ip1(n12321), .ip2(\cache_tag_B[3][18] ), .op(n8175) );
  nand4_1 U8237 ( .ip1(n8178), .ip2(n8177), .ip3(n8176), .ip4(n8175), .op(
        n8179) );
  not_ab_or_c_or_d U8238 ( .ip1(\cache_tag_B[5][18] ), .ip2(n11296), .ip3(
        n8180), .ip4(n8179), .op(n8182) );
  nand2_1 U8239 ( .ip1(n12396), .ip2(\cache_tag_B[4][18] ), .op(n8181) );
  nand3_1 U8240 ( .ip1(n8183), .ip2(n8182), .ip3(n8181), .op(n8184) );
  nand2_1 U8241 ( .ip1(n8545), .ip2(n8184), .op(n8187) );
  nand2_1 U8242 ( .ip1(addr_mem[25]), .ip2(n13201), .op(n8186) );
  nand2_1 U8243 ( .ip1(addr_resp[25]), .ip2(n9703), .op(n8185) );
  nand4_1 U8244 ( .ip1(n8188), .ip2(n8187), .ip3(n8186), .ip4(n8185), .op(
        n5229) );
  nand2_1 U8245 ( .ip1(n12583), .ip2(\cache_tag_B[2][21] ), .op(n8197) );
  inv_1 U8246 ( .ip(\cache_tag_B[7][21] ), .op(n9270) );
  nor2_1 U8247 ( .ip1(n9769), .ip2(n9270), .op(n8194) );
  nand2_1 U8248 ( .ip1(n12321), .ip2(\cache_tag_B[3][21] ), .op(n8192) );
  nand2_1 U8249 ( .ip1(n10686), .ip2(\cache_tag_B[1][21] ), .op(n8191) );
  nand2_1 U8250 ( .ip1(n12256), .ip2(\cache_tag_B[5][21] ), .op(n8190) );
  nand2_1 U8251 ( .ip1(n12396), .ip2(\cache_tag_B[4][21] ), .op(n8189) );
  nand4_1 U8252 ( .ip1(n8192), .ip2(n8191), .ip3(n8190), .ip4(n8189), .op(
        n8193) );
  not_ab_or_c_or_d U8253 ( .ip1(\cache_tag_B[0][21] ), .ip2(n12357), .ip3(
        n8194), .ip4(n8193), .op(n8196) );
  nand2_1 U8254 ( .ip1(n12371), .ip2(\cache_tag_B[6][21] ), .op(n8195) );
  nand3_1 U8255 ( .ip1(n8197), .ip2(n8196), .ip3(n8195), .op(n8198) );
  nand2_1 U8256 ( .ip1(n8545), .ip2(n8198), .op(n8211) );
  nand2_1 U8257 ( .ip1(\cache_tag_A[0][21] ), .ip2(n12204), .op(n8207) );
  inv_1 U8258 ( .ip(\cache_tag_A[6][21] ), .op(n8863) );
  nor2_1 U8259 ( .ip1(n8863), .ip2(n9762), .op(n8204) );
  nand2_1 U8260 ( .ip1(\cache_tag_A[3][21] ), .ip2(n12410), .op(n8202) );
  nand2_1 U8261 ( .ip1(\cache_tag_A[4][21] ), .ip2(n12194), .op(n8201) );
  nand2_1 U8262 ( .ip1(\cache_tag_A[1][21] ), .ip2(n12147), .op(n8200) );
  nand2_1 U8263 ( .ip1(\cache_tag_A[5][21] ), .ip2(n11280), .op(n8199) );
  nand4_1 U8264 ( .ip1(n8202), .ip2(n8201), .ip3(n8200), .ip4(n8199), .op(
        n8203) );
  not_ab_or_c_or_d U8265 ( .ip1(n12278), .ip2(\cache_tag_A[7][21] ), .ip3(
        n8204), .ip4(n8203), .op(n8206) );
  nand2_1 U8266 ( .ip1(\cache_tag_A[2][21] ), .ip2(n12486), .op(n8205) );
  nand3_1 U8267 ( .ip1(n8207), .ip2(n8206), .ip3(n8205), .op(n9462) );
  nand2_1 U8268 ( .ip1(n8555), .ip2(n9462), .op(n8210) );
  nand2_1 U8269 ( .ip1(addr_mem[28]), .ip2(n13201), .op(n8209) );
  nand2_1 U8270 ( .ip1(addr_resp[28]), .ip2(n9619), .op(n8208) );
  nand4_1 U8271 ( .ip1(n8211), .ip2(n8210), .ip3(n8209), .ip4(n8208), .op(
        n5226) );
  nand2_1 U8272 ( .ip1(\cache_tag_A[3][3] ), .ip2(n12410), .op(n8220) );
  inv_1 U8273 ( .ip(n12429), .op(n9762) );
  inv_1 U8274 ( .ip(\cache_tag_A[6][3] ), .op(n8731) );
  nor2_1 U8275 ( .ip1(n9762), .ip2(n8731), .op(n8217) );
  nand2_1 U8276 ( .ip1(n11324), .ip2(\cache_tag_A[4][3] ), .op(n8215) );
  nand2_1 U8277 ( .ip1(n11304), .ip2(\cache_tag_A[5][3] ), .op(n8214) );
  nand2_1 U8278 ( .ip1(n10702), .ip2(\cache_tag_A[7][3] ), .op(n8213) );
  nand2_1 U8279 ( .ip1(n12583), .ip2(\cache_tag_A[2][3] ), .op(n8212) );
  nand4_1 U8280 ( .ip1(n8215), .ip2(n8214), .ip3(n8213), .ip4(n8212), .op(
        n8216) );
  not_ab_or_c_or_d U8281 ( .ip1(\cache_tag_A[0][3] ), .ip2(n12357), .ip3(n8217), .ip4(n8216), .op(n8219) );
  nand2_1 U8282 ( .ip1(n10166), .ip2(\cache_tag_A[1][3] ), .op(n8218) );
  nand3_1 U8283 ( .ip1(n8220), .ip2(n8219), .ip3(n8218), .op(n9512) );
  nand2_1 U8284 ( .ip1(n8555), .ip2(n9512), .op(n8234) );
  nand2_1 U8285 ( .ip1(n12583), .ip2(\cache_tag_B[2][3] ), .op(n8229) );
  inv_1 U8286 ( .ip(\cache_tag_B[7][3] ), .op(n8995) );
  nor2_1 U8287 ( .ip1(n9769), .ip2(n8995), .op(n8226) );
  nand2_1 U8288 ( .ip1(n11946), .ip2(\cache_tag_B[1][3] ), .op(n8224) );
  nand2_1 U8289 ( .ip1(n12584), .ip2(\cache_tag_B[4][3] ), .op(n8223) );
  nand2_1 U8290 ( .ip1(n8452), .ip2(\cache_tag_B[0][3] ), .op(n8222) );
  nand2_1 U8291 ( .ip1(n12591), .ip2(\cache_tag_B[3][3] ), .op(n8221) );
  nand4_1 U8292 ( .ip1(n8224), .ip2(n8223), .ip3(n8222), .ip4(n8221), .op(
        n8225) );
  not_ab_or_c_or_d U8293 ( .ip1(\cache_tag_B[5][3] ), .ip2(n11236), .ip3(n8226), .ip4(n8225), .op(n8228) );
  nand2_1 U8294 ( .ip1(n12551), .ip2(\cache_tag_B[6][3] ), .op(n8227) );
  nand3_1 U8295 ( .ip1(n8229), .ip2(n8228), .ip3(n8227), .op(n8230) );
  nand2_1 U8296 ( .ip1(n8545), .ip2(n8230), .op(n8233) );
  nand2_1 U8297 ( .ip1(addr_mem[10]), .ip2(n13201), .op(n8232) );
  nand2_1 U8298 ( .ip1(addr_resp[10]), .ip2(n9619), .op(n8231) );
  nand4_1 U8299 ( .ip1(n8234), .ip2(n8233), .ip3(n8232), .ip4(n8231), .op(
        n5244) );
  nand2_1 U8300 ( .ip1(n10426), .ip2(\cache_tag_A[2][0] ), .op(n8243) );
  inv_1 U8301 ( .ip(\cache_tag_A[1][0] ), .op(n8742) );
  nor2_1 U8302 ( .ip1(n9862), .ip2(n8742), .op(n8240) );
  nand2_1 U8303 ( .ip1(n11535), .ip2(\cache_tag_A[3][0] ), .op(n8238) );
  buf_1 U8304 ( .ip(n11296), .op(n11280) );
  nand2_1 U8305 ( .ip1(n11280), .ip2(\cache_tag_A[5][0] ), .op(n8237) );
  nand2_1 U8306 ( .ip1(n12458), .ip2(\cache_tag_A[6][0] ), .op(n8236) );
  nand2_1 U8307 ( .ip1(n12370), .ip2(\cache_tag_A[0][0] ), .op(n8235) );
  nand4_1 U8308 ( .ip1(n8238), .ip2(n8237), .ip3(n8236), .ip4(n8235), .op(
        n8239) );
  not_ab_or_c_or_d U8309 ( .ip1(n12278), .ip2(\cache_tag_A[7][0] ), .ip3(n8240), .ip4(n8239), .op(n8242) );
  nand2_1 U8310 ( .ip1(n11324), .ip2(\cache_tag_A[4][0] ), .op(n8241) );
  nand3_1 U8311 ( .ip1(n8243), .ip2(n8242), .ip3(n8241), .op(n9530) );
  nand2_1 U8312 ( .ip1(n8555), .ip2(n9530), .op(n8257) );
  nand2_1 U8313 ( .ip1(n8452), .ip2(\cache_tag_B[0][0] ), .op(n8252) );
  inv_1 U8314 ( .ip(\cache_tag_B[7][0] ), .op(n9076) );
  nor2_1 U8315 ( .ip1(n9769), .ip2(n9076), .op(n8249) );
  nand2_1 U8316 ( .ip1(n12591), .ip2(\cache_tag_B[3][0] ), .op(n8247) );
  nand2_1 U8317 ( .ip1(n11946), .ip2(\cache_tag_B[1][0] ), .op(n8246) );
  nand2_1 U8318 ( .ip1(n12583), .ip2(\cache_tag_B[2][0] ), .op(n8245) );
  nand2_1 U8319 ( .ip1(n12584), .ip2(\cache_tag_B[4][0] ), .op(n8244) );
  nand4_1 U8320 ( .ip1(n8247), .ip2(n8246), .ip3(n8245), .ip4(n8244), .op(
        n8248) );
  not_ab_or_c_or_d U8321 ( .ip1(\cache_tag_B[5][0] ), .ip2(n11236), .ip3(n8249), .ip4(n8248), .op(n8251) );
  nand2_1 U8322 ( .ip1(n12551), .ip2(\cache_tag_B[6][0] ), .op(n8250) );
  nand3_1 U8323 ( .ip1(n8252), .ip2(n8251), .ip3(n8250), .op(n8253) );
  nand2_1 U8324 ( .ip1(n8545), .ip2(n8253), .op(n8256) );
  nand2_1 U8325 ( .ip1(addr_mem[7]), .ip2(n13201), .op(n8255) );
  nand2_1 U8326 ( .ip1(addr_resp[7]), .ip2(n9619), .op(n8254) );
  nand4_1 U8327 ( .ip1(n8257), .ip2(n8256), .ip3(n8255), .ip4(n8254), .op(
        n5247) );
  nand2_1 U8328 ( .ip1(n10166), .ip2(\cache_tag_A[1][1] ), .op(n8266) );
  inv_1 U8329 ( .ip(\cache_tag_A[3][1] ), .op(n8677) );
  nor2_1 U8330 ( .ip1(n9866), .ip2(n8677), .op(n8263) );
  nand2_1 U8331 ( .ip1(n8452), .ip2(\cache_tag_A[0][1] ), .op(n8261) );
  nand2_1 U8332 ( .ip1(n11324), .ip2(\cache_tag_A[4][1] ), .op(n8260) );
  nand2_1 U8333 ( .ip1(n12583), .ip2(\cache_tag_A[2][1] ), .op(n8259) );
  nand2_1 U8334 ( .ip1(n11057), .ip2(\cache_tag_A[7][1] ), .op(n8258) );
  nand4_1 U8335 ( .ip1(n8261), .ip2(n8260), .ip3(n8259), .ip4(n8258), .op(
        n8262) );
  not_ab_or_c_or_d U8336 ( .ip1(\cache_tag_A[6][1] ), .ip2(n12320), .ip3(n8263), .ip4(n8262), .op(n8265) );
  nand2_1 U8337 ( .ip1(n11304), .ip2(\cache_tag_A[5][1] ), .op(n8264) );
  nand3_1 U8338 ( .ip1(n8266), .ip2(n8265), .ip3(n8264), .op(n9492) );
  nand2_1 U8339 ( .ip1(n8555), .ip2(n9492), .op(n8280) );
  nand2_1 U8340 ( .ip1(n12583), .ip2(\cache_tag_B[2][1] ), .op(n8275) );
  inv_1 U8341 ( .ip(\cache_tag_B[7][1] ), .op(n9151) );
  nor2_1 U8342 ( .ip1(n9769), .ip2(n9151), .op(n8272) );
  nand2_1 U8343 ( .ip1(n10686), .ip2(\cache_tag_B[1][1] ), .op(n8270) );
  nand2_1 U8344 ( .ip1(n12357), .ip2(\cache_tag_B[0][1] ), .op(n8269) );
  nand2_1 U8345 ( .ip1(n12584), .ip2(\cache_tag_B[4][1] ), .op(n8268) );
  nand2_1 U8346 ( .ip1(n12591), .ip2(\cache_tag_B[3][1] ), .op(n8267) );
  nand4_1 U8347 ( .ip1(n8270), .ip2(n8269), .ip3(n8268), .ip4(n8267), .op(
        n8271) );
  not_ab_or_c_or_d U8348 ( .ip1(\cache_tag_B[5][1] ), .ip2(n11236), .ip3(n8272), .ip4(n8271), .op(n8274) );
  nand2_1 U8349 ( .ip1(n12551), .ip2(\cache_tag_B[6][1] ), .op(n8273) );
  nand3_1 U8350 ( .ip1(n8275), .ip2(n8274), .ip3(n8273), .op(n8276) );
  nand2_1 U8351 ( .ip1(n8545), .ip2(n8276), .op(n8279) );
  nand2_1 U8352 ( .ip1(addr_mem[8]), .ip2(n13201), .op(n8278) );
  nand2_1 U8353 ( .ip1(addr_resp[8]), .ip2(n9703), .op(n8277) );
  nand4_1 U8354 ( .ip1(n8280), .ip2(n8279), .ip3(n8278), .ip4(n8277), .op(
        n5246) );
  nand2_1 U8355 ( .ip1(n11324), .ip2(\cache_tag_A[4][23] ), .op(n8289) );
  inv_1 U8356 ( .ip(\cache_tag_A[7][23] ), .op(n8949) );
  nor2_1 U8357 ( .ip1(n9769), .ip2(n8949), .op(n8286) );
  nand2_1 U8358 ( .ip1(n12321), .ip2(\cache_tag_A[3][23] ), .op(n8284) );
  nand2_1 U8359 ( .ip1(n12371), .ip2(\cache_tag_A[6][23] ), .op(n8283) );
  nand2_1 U8360 ( .ip1(n12583), .ip2(\cache_tag_A[2][23] ), .op(n8282) );
  nand2_1 U8361 ( .ip1(n11304), .ip2(\cache_tag_A[5][23] ), .op(n8281) );
  nand4_1 U8362 ( .ip1(n8284), .ip2(n8283), .ip3(n8282), .ip4(n8281), .op(
        n8285) );
  not_ab_or_c_or_d U8363 ( .ip1(n12297), .ip2(\cache_tag_A[0][23] ), .ip3(
        n8286), .ip4(n8285), .op(n8288) );
  nand2_1 U8364 ( .ip1(n10166), .ip2(\cache_tag_A[1][23] ), .op(n8287) );
  nand3_1 U8365 ( .ip1(n8289), .ip2(n8288), .ip3(n8287), .op(n9476) );
  nand2_1 U8366 ( .ip1(n8555), .ip2(n9476), .op(n8303) );
  nand2_1 U8367 ( .ip1(n11057), .ip2(\cache_tag_B[7][23] ), .op(n8298) );
  inv_1 U8368 ( .ip(\cache_tag_B[3][23] ), .op(n9242) );
  nor2_1 U8369 ( .ip1(n9866), .ip2(n9242), .op(n8295) );
  nand2_1 U8370 ( .ip1(n11324), .ip2(\cache_tag_B[4][23] ), .op(n8293) );
  nand2_1 U8371 ( .ip1(n12256), .ip2(\cache_tag_B[5][23] ), .op(n8292) );
  nand2_1 U8372 ( .ip1(n12371), .ip2(\cache_tag_B[6][23] ), .op(n8291) );
  nand2_1 U8373 ( .ip1(n12583), .ip2(\cache_tag_B[2][23] ), .op(n8290) );
  nand4_1 U8374 ( .ip1(n8293), .ip2(n8292), .ip3(n8291), .ip4(n8290), .op(
        n8294) );
  not_ab_or_c_or_d U8375 ( .ip1(\cache_tag_B[0][23] ), .ip2(n12357), .ip3(
        n8295), .ip4(n8294), .op(n8297) );
  nand2_1 U8376 ( .ip1(n10166), .ip2(\cache_tag_B[1][23] ), .op(n8296) );
  nand3_1 U8377 ( .ip1(n8298), .ip2(n8297), .ip3(n8296), .op(n8299) );
  nand2_1 U8378 ( .ip1(n8545), .ip2(n8299), .op(n8302) );
  nand2_1 U8379 ( .ip1(addr_mem[30]), .ip2(n13201), .op(n8301) );
  nand2_1 U8380 ( .ip1(addr_resp[30]), .ip2(n9703), .op(n8300) );
  nand4_1 U8381 ( .ip1(n8303), .ip2(n8302), .ip3(n8301), .ip4(n8300), .op(
        n5224) );
  inv_1 U8382 ( .ip(n9769), .op(n12581) );
  buf_1 U8383 ( .ip(n12581), .op(n12468) );
  nand2_1 U8384 ( .ip1(\cache_tag_A[7][12] ), .ip2(n12468), .op(n8312) );
  inv_1 U8385 ( .ip(\cache_tag_A[4][12] ), .op(n8754) );
  nor2_1 U8386 ( .ip1(n9868), .ip2(n8754), .op(n8309) );
  nand2_1 U8387 ( .ip1(n11304), .ip2(\cache_tag_A[5][12] ), .op(n8307) );
  nand2_1 U8388 ( .ip1(n12583), .ip2(\cache_tag_A[2][12] ), .op(n8306) );
  nand2_1 U8389 ( .ip1(n12370), .ip2(\cache_tag_A[0][12] ), .op(n8305) );
  nand2_1 U8390 ( .ip1(n12321), .ip2(\cache_tag_A[3][12] ), .op(n8304) );
  nand4_1 U8391 ( .ip1(n8307), .ip2(n8306), .ip3(n8305), .ip4(n8304), .op(
        n8308) );
  not_ab_or_c_or_d U8392 ( .ip1(n11946), .ip2(\cache_tag_A[1][12] ), .ip3(
        n8309), .ip4(n8308), .op(n8311) );
  nand2_1 U8393 ( .ip1(n12371), .ip2(\cache_tag_A[6][12] ), .op(n8310) );
  nand3_1 U8394 ( .ip1(n8312), .ip2(n8311), .ip3(n8310), .op(n9478) );
  nand2_1 U8395 ( .ip1(n8555), .ip2(n9478), .op(n8326) );
  nand2_1 U8396 ( .ip1(n12194), .ip2(\cache_tag_B[4][12] ), .op(n8321) );
  inv_1 U8397 ( .ip(\cache_tag_B[7][12] ), .op(n9177) );
  nor2_1 U8398 ( .ip1(n9769), .ip2(n9177), .op(n8318) );
  nand2_1 U8399 ( .ip1(n12551), .ip2(\cache_tag_B[6][12] ), .op(n8316) );
  nand2_1 U8400 ( .ip1(n12583), .ip2(\cache_tag_B[2][12] ), .op(n8315) );
  nand2_1 U8401 ( .ip1(n10686), .ip2(\cache_tag_B[1][12] ), .op(n8314) );
  nand2_1 U8402 ( .ip1(n12370), .ip2(\cache_tag_B[0][12] ), .op(n8313) );
  nand4_1 U8403 ( .ip1(n8316), .ip2(n8315), .ip3(n8314), .ip4(n8313), .op(
        n8317) );
  not_ab_or_c_or_d U8404 ( .ip1(\cache_tag_B[3][12] ), .ip2(n12096), .ip3(
        n8318), .ip4(n8317), .op(n8320) );
  nand2_1 U8405 ( .ip1(n12256), .ip2(\cache_tag_B[5][12] ), .op(n8319) );
  nand3_1 U8406 ( .ip1(n8321), .ip2(n8320), .ip3(n8319), .op(n8322) );
  nand2_1 U8407 ( .ip1(n8545), .ip2(n8322), .op(n8325) );
  nand2_1 U8408 ( .ip1(addr_mem[19]), .ip2(n13201), .op(n8324) );
  nand2_1 U8409 ( .ip1(addr_resp[19]), .ip2(n9703), .op(n8323) );
  nand4_1 U8410 ( .ip1(n8326), .ip2(n8325), .ip3(n8324), .ip4(n8323), .op(
        n5235) );
  nand2_1 U8411 ( .ip1(\cache_tag_A[7][17] ), .ip2(n12468), .op(n8335) );
  inv_1 U8412 ( .ip(\cache_tag_A[4][17] ), .op(n8889) );
  nor2_1 U8413 ( .ip1(n9868), .ip2(n8889), .op(n8332) );
  nand2_1 U8414 ( .ip1(n10166), .ip2(\cache_tag_A[1][17] ), .op(n8330) );
  nand2_1 U8415 ( .ip1(n12118), .ip2(\cache_tag_A[5][17] ), .op(n8329) );
  buf_1 U8416 ( .ip(n12370), .op(n11071) );
  nand2_1 U8417 ( .ip1(n11071), .ip2(\cache_tag_A[0][17] ), .op(n8328) );
  nand2_1 U8418 ( .ip1(n12583), .ip2(\cache_tag_A[2][17] ), .op(n8327) );
  nand4_1 U8419 ( .ip1(n8330), .ip2(n8329), .ip3(n8328), .ip4(n8327), .op(
        n8331) );
  not_ab_or_c_or_d U8420 ( .ip1(n12096), .ip2(\cache_tag_A[3][17] ), .ip3(
        n8332), .ip4(n8331), .op(n8334) );
  buf_1 U8421 ( .ip(n12429), .op(n12337) );
  nand2_1 U8422 ( .ip1(n12337), .ip2(\cache_tag_A[6][17] ), .op(n8333) );
  nand3_1 U8423 ( .ip1(n8335), .ip2(n8334), .ip3(n8333), .op(n9468) );
  nand2_1 U8424 ( .ip1(n8555), .ip2(n9468), .op(n8349) );
  nand2_1 U8425 ( .ip1(n12370), .ip2(\cache_tag_B[0][17] ), .op(n8344) );
  inv_1 U8426 ( .ip(\cache_tag_B[7][17] ), .op(n9091) );
  nor2_1 U8427 ( .ip1(n9769), .ip2(n9091), .op(n8341) );
  nand2_1 U8428 ( .ip1(n12256), .ip2(\cache_tag_B[5][17] ), .op(n8339) );
  nand2_1 U8429 ( .ip1(n12551), .ip2(\cache_tag_B[6][17] ), .op(n8338) );
  nand2_1 U8430 ( .ip1(n12396), .ip2(\cache_tag_B[4][17] ), .op(n8337) );
  nand2_1 U8431 ( .ip1(n12321), .ip2(\cache_tag_B[3][17] ), .op(n8336) );
  nand4_1 U8432 ( .ip1(n8339), .ip2(n8338), .ip3(n8337), .ip4(n8336), .op(
        n8340) );
  not_ab_or_c_or_d U8433 ( .ip1(\cache_tag_B[2][17] ), .ip2(n12475), .ip3(
        n8341), .ip4(n8340), .op(n8343) );
  nand2_1 U8434 ( .ip1(n11946), .ip2(\cache_tag_B[1][17] ), .op(n8342) );
  nand3_1 U8435 ( .ip1(n8344), .ip2(n8343), .ip3(n8342), .op(n8345) );
  nand2_1 U8436 ( .ip1(n8545), .ip2(n8345), .op(n8348) );
  nand2_1 U8437 ( .ip1(addr_mem[24]), .ip2(n13201), .op(n8347) );
  nand2_1 U8438 ( .ip1(addr_resp[24]), .ip2(n9703), .op(n8346) );
  nand4_1 U8439 ( .ip1(n8349), .ip2(n8348), .ip3(n8347), .ip4(n8346), .op(
        n5230) );
  nand2_1 U8440 ( .ip1(n12583), .ip2(\cache_tag_B[2][5] ), .op(n8358) );
  inv_1 U8441 ( .ip(\cache_tag_B[5][5] ), .op(n9017) );
  nor2_1 U8442 ( .ip1(n9870), .ip2(n9017), .op(n8355) );
  nand2_1 U8443 ( .ip1(n8452), .ip2(\cache_tag_B[0][5] ), .op(n8353) );
  nand2_1 U8444 ( .ip1(n12584), .ip2(\cache_tag_B[4][5] ), .op(n8352) );
  nand2_1 U8445 ( .ip1(n12591), .ip2(\cache_tag_B[3][5] ), .op(n8351) );
  nand2_1 U8446 ( .ip1(n12551), .ip2(\cache_tag_B[6][5] ), .op(n8350) );
  nand4_1 U8447 ( .ip1(n8353), .ip2(n8352), .ip3(n8351), .ip4(n8350), .op(
        n8354) );
  not_ab_or_c_or_d U8448 ( .ip1(\cache_tag_B[7][5] ), .ip2(n10702), .ip3(n8355), .ip4(n8354), .op(n8357) );
  nand2_1 U8449 ( .ip1(n11946), .ip2(\cache_tag_B[1][5] ), .op(n8356) );
  nand3_1 U8450 ( .ip1(n8358), .ip2(n8357), .ip3(n8356), .op(n8359) );
  nand2_1 U8451 ( .ip1(n8545), .ip2(n8359), .op(n8372) );
  buf_1 U8452 ( .ip(n12581), .op(n12552) );
  nand2_1 U8453 ( .ip1(\cache_tag_A[7][5] ), .ip2(n12552), .op(n8368) );
  inv_1 U8454 ( .ip(\cache_tag_A[5][5] ), .op(n8765) );
  nor2_1 U8455 ( .ip1(n9870), .ip2(n8765), .op(n8365) );
  nand2_1 U8456 ( .ip1(n8452), .ip2(\cache_tag_A[0][5] ), .op(n8363) );
  nand2_1 U8457 ( .ip1(n12583), .ip2(\cache_tag_A[2][5] ), .op(n8362) );
  nand2_1 U8458 ( .ip1(n12371), .ip2(\cache_tag_A[6][5] ), .op(n8361) );
  nand2_1 U8459 ( .ip1(n11324), .ip2(\cache_tag_A[4][5] ), .op(n8360) );
  nand4_1 U8460 ( .ip1(n8363), .ip2(n8362), .ip3(n8361), .ip4(n8360), .op(
        n8364) );
  not_ab_or_c_or_d U8461 ( .ip1(n12096), .ip2(\cache_tag_A[3][5] ), .ip3(n8365), .ip4(n8364), .op(n8367) );
  nand2_1 U8462 ( .ip1(n10166), .ip2(\cache_tag_A[1][5] ), .op(n8366) );
  nand3_1 U8463 ( .ip1(n8368), .ip2(n8367), .ip3(n8366), .op(n9490) );
  nand2_1 U8464 ( .ip1(n8555), .ip2(n9490), .op(n8371) );
  nand2_1 U8465 ( .ip1(addr_mem[12]), .ip2(n13201), .op(n8370) );
  nand2_1 U8466 ( .ip1(addr_resp[12]), .ip2(n9703), .op(n8369) );
  nand4_1 U8467 ( .ip1(n8372), .ip2(n8371), .ip3(n8370), .ip4(n8369), .op(
        n5242) );
  nand2_1 U8468 ( .ip1(\cache_tag_A[7][9] ), .ip2(n12468), .op(n8381) );
  inv_1 U8469 ( .ip(\cache_tag_A[4][9] ), .op(n8814) );
  nor2_1 U8470 ( .ip1(n9868), .ip2(n8814), .op(n8378) );
  nand2_1 U8471 ( .ip1(n8452), .ip2(\cache_tag_A[0][9] ), .op(n8376) );
  nand2_1 U8472 ( .ip1(n11304), .ip2(\cache_tag_A[5][9] ), .op(n8375) );
  nand2_1 U8473 ( .ip1(n12583), .ip2(\cache_tag_A[2][9] ), .op(n8374) );
  nand2_1 U8474 ( .ip1(n10166), .ip2(\cache_tag_A[1][9] ), .op(n8373) );
  nand4_1 U8475 ( .ip1(n8376), .ip2(n8375), .ip3(n8374), .ip4(n8373), .op(
        n8377) );
  not_ab_or_c_or_d U8476 ( .ip1(\cache_tag_A[3][9] ), .ip2(n12096), .ip3(n8378), .ip4(n8377), .op(n8380) );
  nand2_1 U8477 ( .ip1(n12371), .ip2(\cache_tag_A[6][9] ), .op(n8379) );
  nand3_1 U8478 ( .ip1(n8381), .ip2(n8380), .ip3(n8379), .op(n9500) );
  nand2_1 U8479 ( .ip1(n8555), .ip2(n9500), .op(n8395) );
  nand2_1 U8480 ( .ip1(n12591), .ip2(\cache_tag_B[3][9] ), .op(n8390) );
  inv_1 U8481 ( .ip(\cache_tag_B[7][9] ), .op(n9114) );
  nor2_1 U8482 ( .ip1(n9769), .ip2(n9114), .op(n8387) );
  nand2_1 U8483 ( .ip1(n12583), .ip2(\cache_tag_B[2][9] ), .op(n8385) );
  nand2_1 U8484 ( .ip1(n11946), .ip2(\cache_tag_B[1][9] ), .op(n8384) );
  nand2_1 U8485 ( .ip1(n12370), .ip2(\cache_tag_B[0][9] ), .op(n8383) );
  nand2_1 U8486 ( .ip1(n12551), .ip2(\cache_tag_B[6][9] ), .op(n8382) );
  nand4_1 U8487 ( .ip1(n8385), .ip2(n8384), .ip3(n8383), .ip4(n8382), .op(
        n8386) );
  not_ab_or_c_or_d U8488 ( .ip1(\cache_tag_B[4][9] ), .ip2(n12194), .ip3(n8387), .ip4(n8386), .op(n8389) );
  nand2_1 U8489 ( .ip1(n12118), .ip2(\cache_tag_B[5][9] ), .op(n8388) );
  nand3_1 U8490 ( .ip1(n8390), .ip2(n8389), .ip3(n8388), .op(n8391) );
  nand2_1 U8491 ( .ip1(n8545), .ip2(n8391), .op(n8394) );
  nand2_1 U8492 ( .ip1(addr_mem[16]), .ip2(n13201), .op(n8393) );
  nand2_1 U8493 ( .ip1(addr_resp[16]), .ip2(n9703), .op(n8392) );
  nand4_1 U8494 ( .ip1(n8395), .ip2(n8394), .ip3(n8393), .ip4(n8392), .op(
        n5238) );
  nand2_1 U8495 ( .ip1(addr_mem[18]), .ip2(n13201), .op(n8418) );
  nand2_1 U8496 ( .ip1(n11057), .ip2(\cache_tag_A[7][11] ), .op(n8404) );
  inv_1 U8497 ( .ip(\cache_tag_A[6][11] ), .op(n8792) );
  nor2_1 U8498 ( .ip1(n9762), .ip2(n8792), .op(n8401) );
  nand2_1 U8499 ( .ip1(n12410), .ip2(\cache_tag_A[3][11] ), .op(n8399) );
  nand2_1 U8500 ( .ip1(n12583), .ip2(\cache_tag_A[2][11] ), .op(n8398) );
  nand2_1 U8501 ( .ip1(n8452), .ip2(\cache_tag_A[0][11] ), .op(n8397) );
  nand2_1 U8502 ( .ip1(n11304), .ip2(\cache_tag_A[5][11] ), .op(n8396) );
  nand4_1 U8503 ( .ip1(n8399), .ip2(n8398), .ip3(n8397), .ip4(n8396), .op(
        n8400) );
  not_ab_or_c_or_d U8504 ( .ip1(n11946), .ip2(\cache_tag_A[1][11] ), .ip3(
        n8401), .ip4(n8400), .op(n8403) );
  nand2_1 U8505 ( .ip1(n11324), .ip2(\cache_tag_A[4][11] ), .op(n8402) );
  nand3_1 U8506 ( .ip1(n8404), .ip2(n8403), .ip3(n8402), .op(n9488) );
  nand2_1 U8507 ( .ip1(n8555), .ip2(n9488), .op(n8417) );
  nand2_1 U8508 ( .ip1(n12320), .ip2(\cache_tag_B[6][11] ), .op(n8413) );
  inv_1 U8509 ( .ip(\cache_tag_B[7][11] ), .op(n9190) );
  nor2_1 U8510 ( .ip1(n9769), .ip2(n9190), .op(n8410) );
  nand2_1 U8511 ( .ip1(n12591), .ip2(\cache_tag_B[3][11] ), .op(n8408) );
  nand2_1 U8512 ( .ip1(n12370), .ip2(\cache_tag_B[0][11] ), .op(n8407) );
  nand2_1 U8513 ( .ip1(n12583), .ip2(\cache_tag_B[2][11] ), .op(n8406) );
  nand2_1 U8514 ( .ip1(n12256), .ip2(\cache_tag_B[5][11] ), .op(n8405) );
  nand4_1 U8515 ( .ip1(n8408), .ip2(n8407), .ip3(n8406), .ip4(n8405), .op(
        n8409) );
  not_ab_or_c_or_d U8516 ( .ip1(\cache_tag_B[1][11] ), .ip2(n11946), .ip3(
        n8410), .ip4(n8409), .op(n8412) );
  nand2_1 U8517 ( .ip1(n12396), .ip2(\cache_tag_B[4][11] ), .op(n8411) );
  nand3_1 U8518 ( .ip1(n8413), .ip2(n8412), .ip3(n8411), .op(n8414) );
  nand2_1 U8519 ( .ip1(n8545), .ip2(n8414), .op(n8416) );
  nand2_1 U8520 ( .ip1(addr_resp[18]), .ip2(n9703), .op(n8415) );
  nand4_1 U8521 ( .ip1(n8418), .ip2(n8417), .ip3(n8416), .ip4(n8415), .op(
        n5236) );
  nand2_1 U8522 ( .ip1(addr_mem[15]), .ip2(n13201), .op(n8441) );
  nand2_1 U8523 ( .ip1(n12204), .ip2(\cache_tag_A[0][8] ), .op(n8427) );
  inv_1 U8524 ( .ip(\cache_tag_A[6][8] ), .op(n8825) );
  nor2_1 U8525 ( .ip1(n9762), .ip2(n8825), .op(n8424) );
  nand2_1 U8526 ( .ip1(n11304), .ip2(\cache_tag_A[5][8] ), .op(n8422) );
  nand2_1 U8527 ( .ip1(n12054), .ip2(\cache_tag_A[4][8] ), .op(n8421) );
  nand2_1 U8528 ( .ip1(n12321), .ip2(\cache_tag_A[3][8] ), .op(n8420) );
  buf_1 U8529 ( .ip(n11724), .op(n10686) );
  nand2_1 U8530 ( .ip1(n10686), .ip2(\cache_tag_A[1][8] ), .op(n8419) );
  nand4_1 U8531 ( .ip1(n8422), .ip2(n8421), .ip3(n8420), .ip4(n8419), .op(
        n8423) );
  not_ab_or_c_or_d U8532 ( .ip1(\cache_tag_A[7][8] ), .ip2(n11057), .ip3(n8424), .ip4(n8423), .op(n8426) );
  buf_1 U8533 ( .ip(n12546), .op(n11142) );
  nand2_1 U8534 ( .ip1(n11142), .ip2(\cache_tag_A[2][8] ), .op(n8425) );
  nand3_1 U8535 ( .ip1(n8427), .ip2(n8426), .ip3(n8425), .op(n9466) );
  nand2_1 U8536 ( .ip1(n8555), .ip2(n9466), .op(n8440) );
  nand2_1 U8537 ( .ip1(n11780), .ip2(\cache_tag_B[6][8] ), .op(n8436) );
  inv_1 U8538 ( .ip(\cache_tag_B[7][8] ), .op(n9125) );
  nor2_1 U8539 ( .ip1(n9769), .ip2(n9125), .op(n8433) );
  nand2_1 U8540 ( .ip1(n8452), .ip2(\cache_tag_B[0][8] ), .op(n8431) );
  nand2_1 U8541 ( .ip1(n12583), .ip2(\cache_tag_B[2][8] ), .op(n8430) );
  nand2_1 U8542 ( .ip1(n12396), .ip2(\cache_tag_B[4][8] ), .op(n8429) );
  nand2_1 U8543 ( .ip1(n10686), .ip2(\cache_tag_B[1][8] ), .op(n8428) );
  nand4_1 U8544 ( .ip1(n8431), .ip2(n8430), .ip3(n8429), .ip4(n8428), .op(
        n8432) );
  not_ab_or_c_or_d U8545 ( .ip1(\cache_tag_B[5][8] ), .ip2(n11236), .ip3(n8433), .ip4(n8432), .op(n8435) );
  nand2_1 U8546 ( .ip1(n12591), .ip2(\cache_tag_B[3][8] ), .op(n8434) );
  nand3_1 U8547 ( .ip1(n8436), .ip2(n8435), .ip3(n8434), .op(n8437) );
  nand2_1 U8548 ( .ip1(n8545), .ip2(n8437), .op(n8439) );
  nand2_1 U8549 ( .ip1(addr_resp[15]), .ip2(n9703), .op(n8438) );
  nand4_1 U8550 ( .ip1(n8441), .ip2(n8440), .ip3(n8439), .ip4(n8438), .op(
        n5239) );
  nand2_1 U8551 ( .ip1(n12583), .ip2(\cache_tag_B[2][20] ), .op(n8450) );
  inv_1 U8552 ( .ip(\cache_tag_B[7][20] ), .op(n9006) );
  nor2_1 U8553 ( .ip1(n9769), .ip2(n9006), .op(n8447) );
  nand2_1 U8554 ( .ip1(n10686), .ip2(\cache_tag_B[1][20] ), .op(n8445) );
  nand2_1 U8555 ( .ip1(n12370), .ip2(\cache_tag_B[0][20] ), .op(n8444) );
  nand2_1 U8556 ( .ip1(n12396), .ip2(\cache_tag_B[4][20] ), .op(n8443) );
  nand2_1 U8557 ( .ip1(n12256), .ip2(\cache_tag_B[5][20] ), .op(n8442) );
  nand4_1 U8558 ( .ip1(n8445), .ip2(n8444), .ip3(n8443), .ip4(n8442), .op(
        n8446) );
  not_ab_or_c_or_d U8559 ( .ip1(\cache_tag_B[3][20] ), .ip2(n12096), .ip3(
        n8447), .ip4(n8446), .op(n8449) );
  nand2_1 U8560 ( .ip1(n12371), .ip2(\cache_tag_B[6][20] ), .op(n8448) );
  nand3_1 U8561 ( .ip1(n8450), .ip2(n8449), .ip3(n8448), .op(n8451) );
  nand2_1 U8562 ( .ip1(n8545), .ip2(n8451), .op(n8465) );
  nand2_1 U8563 ( .ip1(\cache_tag_A[1][20] ), .ip2(n12147), .op(n8461) );
  nand2_1 U8564 ( .ip1(n11304), .ip2(\cache_tag_A[5][20] ), .op(n8460) );
  inv_1 U8565 ( .ip(\cache_tag_A[4][20] ), .op(n8972) );
  nor2_1 U8566 ( .ip1(n9868), .ip2(n8972), .op(n8458) );
  nand2_1 U8567 ( .ip1(n8452), .ip2(\cache_tag_A[0][20] ), .op(n8456) );
  nand2_1 U8568 ( .ip1(n12371), .ip2(\cache_tag_A[6][20] ), .op(n8455) );
  nand2_1 U8569 ( .ip1(n12583), .ip2(\cache_tag_A[2][20] ), .op(n8454) );
  nand2_1 U8570 ( .ip1(n12410), .ip2(\cache_tag_A[3][20] ), .op(n8453) );
  nand4_1 U8571 ( .ip1(n8456), .ip2(n8455), .ip3(n8454), .ip4(n8453), .op(
        n8457) );
  not_ab_or_c_or_d U8572 ( .ip1(n12278), .ip2(\cache_tag_A[7][20] ), .ip3(
        n8458), .ip4(n8457), .op(n8459) );
  nand3_1 U8573 ( .ip1(n8461), .ip2(n8460), .ip3(n8459), .op(n9494) );
  nand2_1 U8574 ( .ip1(n8555), .ip2(n9494), .op(n8464) );
  nand2_1 U8575 ( .ip1(addr_mem[27]), .ip2(n13201), .op(n8463) );
  nand2_1 U8576 ( .ip1(addr_resp[27]), .ip2(n9703), .op(n8462) );
  nand4_1 U8577 ( .ip1(n8465), .ip2(n8464), .ip3(n8463), .ip4(n8462), .op(
        n5227) );
  nand2_1 U8578 ( .ip1(n12321), .ip2(\cache_tag_A[3][19] ), .op(n8474) );
  inv_1 U8579 ( .ip(\cache_tag_A[1][19] ), .op(n8923) );
  nor2_1 U8580 ( .ip1(n9862), .ip2(n8923), .op(n8471) );
  nand2_1 U8581 ( .ip1(n12370), .ip2(\cache_tag_A[0][19] ), .op(n8469) );
  nand2_1 U8582 ( .ip1(n11324), .ip2(\cache_tag_A[4][19] ), .op(n8468) );
  nand2_1 U8583 ( .ip1(n12583), .ip2(\cache_tag_A[2][19] ), .op(n8467) );
  nand2_1 U8584 ( .ip1(n10575), .ip2(\cache_tag_A[7][19] ), .op(n8466) );
  nand4_1 U8585 ( .ip1(n8469), .ip2(n8468), .ip3(n8467), .ip4(n8466), .op(
        n8470) );
  not_ab_or_c_or_d U8586 ( .ip1(n12551), .ip2(\cache_tag_A[6][19] ), .ip3(
        n8471), .ip4(n8470), .op(n8473) );
  nand2_1 U8587 ( .ip1(n11304), .ip2(\cache_tag_A[5][19] ), .op(n8472) );
  nand3_1 U8588 ( .ip1(n8474), .ip2(n8473), .ip3(n8472), .op(n9480) );
  nand2_1 U8589 ( .ip1(n8555), .ip2(n9480), .op(n8488) );
  nand2_1 U8590 ( .ip1(n12458), .ip2(\cache_tag_B[6][19] ), .op(n8483) );
  inv_1 U8591 ( .ip(\cache_tag_B[7][19] ), .op(n9065) );
  nor2_1 U8592 ( .ip1(n9769), .ip2(n9065), .op(n8480) );
  nand2_1 U8593 ( .ip1(n12396), .ip2(\cache_tag_B[4][19] ), .op(n8478) );
  nand2_1 U8594 ( .ip1(n12370), .ip2(\cache_tag_B[0][19] ), .op(n8477) );
  nand2_1 U8595 ( .ip1(n12321), .ip2(\cache_tag_B[3][19] ), .op(n8476) );
  nand2_1 U8596 ( .ip1(n12583), .ip2(\cache_tag_B[2][19] ), .op(n8475) );
  nand4_1 U8597 ( .ip1(n8478), .ip2(n8477), .ip3(n8476), .ip4(n8475), .op(
        n8479) );
  not_ab_or_c_or_d U8598 ( .ip1(\cache_tag_B[1][19] ), .ip2(n11946), .ip3(
        n8480), .ip4(n8479), .op(n8482) );
  nand2_1 U8599 ( .ip1(n12256), .ip2(\cache_tag_B[5][19] ), .op(n8481) );
  nand3_1 U8600 ( .ip1(n8483), .ip2(n8482), .ip3(n8481), .op(n8484) );
  nand2_1 U8601 ( .ip1(n8545), .ip2(n8484), .op(n8487) );
  nand2_1 U8602 ( .ip1(addr_mem[26]), .ip2(n13201), .op(n8486) );
  nand2_1 U8603 ( .ip1(addr_resp[26]), .ip2(n9703), .op(n8485) );
  nand4_1 U8604 ( .ip1(n8488), .ip2(n8487), .ip3(n8486), .ip4(n8485), .op(
        n5228) );
  nand2_1 U8605 ( .ip1(addr_mem[14]), .ip2(n13201), .op(n8511) );
  nand2_1 U8606 ( .ip1(n10702), .ip2(\cache_tag_B[7][7] ), .op(n8497) );
  and2_1 U8607 ( .ip1(n12486), .ip2(\cache_tag_B[2][7] ), .op(n8494) );
  nand2_1 U8608 ( .ip1(n12591), .ip2(\cache_tag_B[3][7] ), .op(n8492) );
  nand2_1 U8609 ( .ip1(n11946), .ip2(\cache_tag_B[1][7] ), .op(n8491) );
  nand2_1 U8610 ( .ip1(n12396), .ip2(\cache_tag_B[4][7] ), .op(n8490) );
  nand2_1 U8611 ( .ip1(n12370), .ip2(\cache_tag_B[0][7] ), .op(n8489) );
  nand4_1 U8612 ( .ip1(n8492), .ip2(n8491), .ip3(n8490), .ip4(n8489), .op(
        n8493) );
  not_ab_or_c_or_d U8613 ( .ip1(\cache_tag_B[5][7] ), .ip2(n11236), .ip3(n8494), .ip4(n8493), .op(n8496) );
  nand2_1 U8614 ( .ip1(n12458), .ip2(\cache_tag_B[6][7] ), .op(n8495) );
  nand3_1 U8615 ( .ip1(n8497), .ip2(n8496), .ip3(n8495), .op(n8498) );
  nand2_1 U8616 ( .ip1(n8545), .ip2(n8498), .op(n8510) );
  nand2_1 U8617 ( .ip1(\cache_tag_A[0][7] ), .ip2(n12204), .op(n8507) );
  inv_1 U8618 ( .ip(\cache_tag_A[4][7] ), .op(n8851) );
  nor2_1 U8619 ( .ip1(n9868), .ip2(n8851), .op(n8504) );
  nand2_1 U8620 ( .ip1(n12321), .ip2(\cache_tag_A[3][7] ), .op(n8502) );
  nand2_1 U8621 ( .ip1(n11057), .ip2(\cache_tag_A[7][7] ), .op(n8501) );
  nand2_1 U8622 ( .ip1(n12371), .ip2(\cache_tag_A[6][7] ), .op(n8500) );
  nand2_1 U8623 ( .ip1(n10166), .ip2(\cache_tag_A[1][7] ), .op(n8499) );
  nand4_1 U8624 ( .ip1(n8502), .ip2(n8501), .ip3(n8500), .ip4(n8499), .op(
        n8503) );
  not_ab_or_c_or_d U8625 ( .ip1(n12546), .ip2(\cache_tag_A[2][7] ), .ip3(n8504), .ip4(n8503), .op(n8506) );
  nand2_1 U8626 ( .ip1(n11304), .ip2(\cache_tag_A[5][7] ), .op(n8505) );
  nand3_1 U8627 ( .ip1(n8507), .ip2(n8506), .ip3(n8505), .op(n9482) );
  nand2_1 U8628 ( .ip1(n8555), .ip2(n9482), .op(n8509) );
  nand2_1 U8629 ( .ip1(addr_resp[14]), .ip2(n9703), .op(n8508) );
  nand4_1 U8630 ( .ip1(n8511), .ip2(n8510), .ip3(n8509), .ip4(n8508), .op(
        n5240) );
  nand2_1 U8631 ( .ip1(addr_mem[17]), .ip2(n13201), .op(n8534) );
  nand2_1 U8632 ( .ip1(\cache_tag_A[4][10] ), .ip2(n12194), .op(n8520) );
  inv_1 U8633 ( .ip(\cache_tag_A[3][10] ), .op(n8803) );
  nor2_1 U8634 ( .ip1(n9866), .ip2(n8803), .op(n8517) );
  nand2_1 U8635 ( .ip1(n10702), .ip2(\cache_tag_A[7][10] ), .op(n8515) );
  nand2_1 U8636 ( .ip1(n11304), .ip2(\cache_tag_A[5][10] ), .op(n8514) );
  nand2_1 U8637 ( .ip1(n12458), .ip2(\cache_tag_A[6][10] ), .op(n8513) );
  nand2_1 U8638 ( .ip1(n12583), .ip2(\cache_tag_A[2][10] ), .op(n8512) );
  nand4_1 U8639 ( .ip1(n8515), .ip2(n8514), .ip3(n8513), .ip4(n8512), .op(
        n8516) );
  not_ab_or_c_or_d U8640 ( .ip1(\cache_tag_A[0][10] ), .ip2(n12357), .ip3(
        n8517), .ip4(n8516), .op(n8519) );
  nand2_1 U8641 ( .ip1(n10166), .ip2(\cache_tag_A[1][10] ), .op(n8518) );
  nand3_1 U8642 ( .ip1(n8520), .ip2(n8519), .ip3(n8518), .op(n9524) );
  nand2_1 U8643 ( .ip1(n8555), .ip2(n9524), .op(n8533) );
  nand2_1 U8644 ( .ip1(n12591), .ip2(\cache_tag_B[3][10] ), .op(n8529) );
  inv_1 U8645 ( .ip(\cache_tag_B[7][10] ), .op(n9283) );
  nor2_1 U8646 ( .ip1(n9769), .ip2(n9283), .op(n8526) );
  nand2_1 U8647 ( .ip1(n11780), .ip2(\cache_tag_B[6][10] ), .op(n8524) );
  nand2_1 U8648 ( .ip1(n12583), .ip2(\cache_tag_B[2][10] ), .op(n8523) );
  nand2_1 U8649 ( .ip1(n12370), .ip2(\cache_tag_B[0][10] ), .op(n8522) );
  nand2_1 U8650 ( .ip1(n12396), .ip2(\cache_tag_B[4][10] ), .op(n8521) );
  nand4_1 U8651 ( .ip1(n8524), .ip2(n8523), .ip3(n8522), .ip4(n8521), .op(
        n8525) );
  not_ab_or_c_or_d U8652 ( .ip1(\cache_tag_B[1][10] ), .ip2(n11946), .ip3(
        n8526), .ip4(n8525), .op(n8528) );
  nand2_1 U8653 ( .ip1(n12256), .ip2(\cache_tag_B[5][10] ), .op(n8527) );
  nand3_1 U8654 ( .ip1(n8529), .ip2(n8528), .ip3(n8527), .op(n8530) );
  nand2_1 U8655 ( .ip1(n8545), .ip2(n8530), .op(n8532) );
  nand2_1 U8656 ( .ip1(addr_resp[17]), .ip2(n9703), .op(n8531) );
  nand4_1 U8657 ( .ip1(n8534), .ip2(n8533), .ip3(n8532), .ip4(n8531), .op(
        n5237) );
  nand2_1 U8658 ( .ip1(n12591), .ip2(\cache_tag_B[3][13] ), .op(n8543) );
  inv_1 U8659 ( .ip(\cache_tag_B[7][13] ), .op(n9258) );
  nor2_1 U8660 ( .ip1(n9769), .ip2(n9258), .op(n8540) );
  nand2_1 U8661 ( .ip1(n12320), .ip2(\cache_tag_B[6][13] ), .op(n8538) );
  nand2_1 U8662 ( .ip1(n12396), .ip2(\cache_tag_B[4][13] ), .op(n8537) );
  nand2_1 U8663 ( .ip1(n12583), .ip2(\cache_tag_B[2][13] ), .op(n8536) );
  nand2_1 U8664 ( .ip1(n12370), .ip2(\cache_tag_B[0][13] ), .op(n8535) );
  nand4_1 U8665 ( .ip1(n8538), .ip2(n8537), .ip3(n8536), .ip4(n8535), .op(
        n8539) );
  not_ab_or_c_or_d U8666 ( .ip1(\cache_tag_B[5][13] ), .ip2(n11296), .ip3(
        n8540), .ip4(n8539), .op(n8542) );
  nand2_1 U8667 ( .ip1(n10686), .ip2(\cache_tag_B[1][13] ), .op(n8541) );
  nand3_1 U8668 ( .ip1(n8543), .ip2(n8542), .ip3(n8541), .op(n8544) );
  nand2_1 U8669 ( .ip1(n8545), .ip2(n8544), .op(n8559) );
  nand2_1 U8670 ( .ip1(n12370), .ip2(\cache_tag_A[0][13] ), .op(n8554) );
  inv_1 U8671 ( .ip(\cache_tag_A[5][13] ), .op(n8911) );
  nor2_1 U8672 ( .ip1(n9870), .ip2(n8911), .op(n8551) );
  nand2_1 U8673 ( .ip1(n10702), .ip2(\cache_tag_A[7][13] ), .op(n8549) );
  nand2_1 U8674 ( .ip1(n11324), .ip2(\cache_tag_A[4][13] ), .op(n8548) );
  nand2_1 U8675 ( .ip1(n11535), .ip2(\cache_tag_A[3][13] ), .op(n8547) );
  nand2_1 U8676 ( .ip1(n11724), .ip2(\cache_tag_A[1][13] ), .op(n8546) );
  nand4_1 U8677 ( .ip1(n8549), .ip2(n8548), .ip3(n8547), .ip4(n8546), .op(
        n8550) );
  not_ab_or_c_or_d U8678 ( .ip1(\cache_tag_A[6][13] ), .ip2(n12320), .ip3(
        n8551), .ip4(n8550), .op(n8553) );
  nand2_1 U8679 ( .ip1(n12583), .ip2(\cache_tag_A[2][13] ), .op(n8552) );
  nand3_1 U8680 ( .ip1(n8554), .ip2(n8553), .ip3(n8552), .op(n9516) );
  nand2_1 U8681 ( .ip1(n8555), .ip2(n9516), .op(n8558) );
  nand2_1 U8682 ( .ip1(addr_mem[20]), .ip2(n13201), .op(n8557) );
  nand2_1 U8683 ( .ip1(addr_resp[20]), .ip2(n9703), .op(n8556) );
  nand4_1 U8684 ( .ip1(n8559), .ip2(n8558), .ip3(n8557), .ip4(n8556), .op(
        n5234) );
  buf_1 U8685 ( .ip(n13297), .op(n13298) );
  buf_1 U8686 ( .ip(rst), .op(n13296) );
  buf_1 U8687 ( .ip(rst), .op(n13297) );
  nand2_1 U8688 ( .ip1(n8620), .ip2(hit), .op(n8560) );
  and3_1 U8689 ( .ip1(n8620), .ip2(hit), .ip3(cache_hit_count[0]), .op(n13250)
         );
  or2_1 U8690 ( .ip1(n8560), .ip2(n13250), .op(n8563) );
  inv_1 U8691 ( .ip(cache_hit_count[0]), .op(n8561) );
  or2_1 U8692 ( .ip1(n8561), .ip2(n13250), .op(n8562) );
  nand2_1 U8693 ( .ip1(n8563), .ip2(n8562), .op(n5156) );
  nand2_1 U8694 ( .ip1(n13250), .ip2(cache_hit_count[1]), .op(n8564) );
  inv_1 U8695 ( .ip(cache_hit_count[2]), .op(n8565) );
  nor2_1 U8696 ( .ip1(n8564), .ip2(n8565), .op(n13249) );
  or2_1 U8697 ( .ip1(n8564), .ip2(n13249), .op(n8567) );
  or2_1 U8698 ( .ip1(n8565), .ip2(n13249), .op(n8566) );
  nand2_1 U8699 ( .ip1(n8567), .ip2(n8566), .op(n5158) );
  nand2_1 U8700 ( .ip1(n13249), .ip2(cache_hit_count[3]), .op(n8568) );
  inv_1 U8701 ( .ip(cache_hit_count[4]), .op(n8569) );
  nor2_1 U8702 ( .ip1(n8568), .ip2(n8569), .op(n13248) );
  or2_1 U8703 ( .ip1(n8568), .ip2(n13248), .op(n8571) );
  or2_1 U8704 ( .ip1(n8569), .ip2(n13248), .op(n8570) );
  nand2_1 U8705 ( .ip1(n8571), .ip2(n8570), .op(n5160) );
  nand2_1 U8706 ( .ip1(n13248), .ip2(cache_hit_count[5]), .op(n8572) );
  inv_1 U8707 ( .ip(cache_hit_count[6]), .op(n8573) );
  nor2_1 U8708 ( .ip1(n8572), .ip2(n8573), .op(n13247) );
  or2_1 U8709 ( .ip1(n8572), .ip2(n13247), .op(n8575) );
  or2_1 U8710 ( .ip1(n8573), .ip2(n13247), .op(n8574) );
  nand2_1 U8711 ( .ip1(n8575), .ip2(n8574), .op(n5162) );
  nand2_1 U8712 ( .ip1(n13247), .ip2(cache_hit_count[7]), .op(n8576) );
  inv_1 U8713 ( .ip(cache_hit_count[8]), .op(n8577) );
  nor2_1 U8714 ( .ip1(n8576), .ip2(n8577), .op(n13246) );
  or2_1 U8715 ( .ip1(n8576), .ip2(n13246), .op(n8579) );
  or2_1 U8716 ( .ip1(n8577), .ip2(n13246), .op(n8578) );
  nand2_1 U8717 ( .ip1(n8579), .ip2(n8578), .op(n5164) );
  nand2_1 U8718 ( .ip1(n13246), .ip2(cache_hit_count[9]), .op(n8580) );
  inv_1 U8719 ( .ip(cache_hit_count[10]), .op(n8581) );
  nor2_1 U8720 ( .ip1(n8580), .ip2(n8581), .op(n13245) );
  or2_1 U8721 ( .ip1(n8580), .ip2(n13245), .op(n8583) );
  or2_1 U8722 ( .ip1(n8581), .ip2(n13245), .op(n8582) );
  nand2_1 U8723 ( .ip1(n8583), .ip2(n8582), .op(n5166) );
  nand2_1 U8724 ( .ip1(n13245), .ip2(cache_hit_count[11]), .op(n8584) );
  inv_1 U8725 ( .ip(cache_hit_count[12]), .op(n8585) );
  nor2_1 U8726 ( .ip1(n8584), .ip2(n8585), .op(n13244) );
  or2_1 U8727 ( .ip1(n8584), .ip2(n13244), .op(n8587) );
  or2_1 U8728 ( .ip1(n8585), .ip2(n13244), .op(n8586) );
  nand2_1 U8729 ( .ip1(n8587), .ip2(n8586), .op(n5168) );
  nand2_1 U8730 ( .ip1(n13244), .ip2(cache_hit_count[13]), .op(n8588) );
  inv_1 U8731 ( .ip(cache_hit_count[14]), .op(n8589) );
  nor2_1 U8732 ( .ip1(n8588), .ip2(n8589), .op(n13243) );
  or2_1 U8733 ( .ip1(n8588), .ip2(n13243), .op(n8591) );
  or2_1 U8734 ( .ip1(n8589), .ip2(n13243), .op(n8590) );
  nand2_1 U8735 ( .ip1(n8591), .ip2(n8590), .op(n5170) );
  nand2_1 U8736 ( .ip1(n13243), .ip2(cache_hit_count[15]), .op(n8592) );
  inv_1 U8737 ( .ip(cache_hit_count[16]), .op(n8593) );
  nor2_1 U8738 ( .ip1(n8592), .ip2(n8593), .op(n13242) );
  or2_1 U8739 ( .ip1(n8592), .ip2(n13242), .op(n8595) );
  or2_1 U8740 ( .ip1(n8593), .ip2(n13242), .op(n8594) );
  nand2_1 U8741 ( .ip1(n8595), .ip2(n8594), .op(n5172) );
  nand2_1 U8742 ( .ip1(n13242), .ip2(cache_hit_count[17]), .op(n8596) );
  inv_1 U8743 ( .ip(cache_hit_count[18]), .op(n8597) );
  nor2_1 U8744 ( .ip1(n8596), .ip2(n8597), .op(n13241) );
  or2_1 U8745 ( .ip1(n8596), .ip2(n13241), .op(n8599) );
  or2_1 U8746 ( .ip1(n8597), .ip2(n13241), .op(n8598) );
  nand2_1 U8747 ( .ip1(n8599), .ip2(n8598), .op(n5174) );
  nand2_1 U8748 ( .ip1(n13241), .ip2(cache_hit_count[19]), .op(n8600) );
  inv_1 U8749 ( .ip(cache_hit_count[20]), .op(n8601) );
  nor2_1 U8750 ( .ip1(n8600), .ip2(n8601), .op(n13240) );
  or2_1 U8751 ( .ip1(n8600), .ip2(n13240), .op(n8603) );
  or2_1 U8752 ( .ip1(n8601), .ip2(n13240), .op(n8602) );
  nand2_1 U8753 ( .ip1(n8603), .ip2(n8602), .op(n5176) );
  nand2_1 U8754 ( .ip1(n13240), .ip2(cache_hit_count[21]), .op(n8604) );
  inv_1 U8755 ( .ip(cache_hit_count[22]), .op(n8605) );
  nor2_1 U8756 ( .ip1(n8604), .ip2(n8605), .op(n13239) );
  or2_1 U8757 ( .ip1(n8604), .ip2(n13239), .op(n8607) );
  or2_1 U8758 ( .ip1(n8605), .ip2(n13239), .op(n8606) );
  nand2_1 U8759 ( .ip1(n8607), .ip2(n8606), .op(n5178) );
  nand2_1 U8760 ( .ip1(n13239), .ip2(cache_hit_count[23]), .op(n8608) );
  inv_1 U8761 ( .ip(cache_hit_count[24]), .op(n8609) );
  nor2_1 U8762 ( .ip1(n8608), .ip2(n8609), .op(n13238) );
  or2_1 U8763 ( .ip1(n8608), .ip2(n13238), .op(n8611) );
  or2_1 U8764 ( .ip1(n8609), .ip2(n13238), .op(n8610) );
  nand2_1 U8765 ( .ip1(n8611), .ip2(n8610), .op(n5180) );
  nand2_1 U8766 ( .ip1(n13238), .ip2(cache_hit_count[25]), .op(n8612) );
  inv_1 U8767 ( .ip(cache_hit_count[26]), .op(n8613) );
  nor2_1 U8768 ( .ip1(n8612), .ip2(n8613), .op(n13237) );
  or2_1 U8769 ( .ip1(n8612), .ip2(n13237), .op(n8615) );
  or2_1 U8770 ( .ip1(n8613), .ip2(n13237), .op(n8614) );
  nand2_1 U8771 ( .ip1(n8615), .ip2(n8614), .op(n5182) );
  nand2_1 U8772 ( .ip1(n13237), .ip2(cache_hit_count[27]), .op(n8616) );
  inv_1 U8773 ( .ip(cache_hit_count[28]), .op(n8617) );
  nor2_1 U8774 ( .ip1(n8616), .ip2(n8617), .op(n13236) );
  or2_1 U8775 ( .ip1(n8616), .ip2(n13236), .op(n8619) );
  or2_1 U8776 ( .ip1(n8617), .ip2(n13236), .op(n8618) );
  nand2_1 U8777 ( .ip1(n8619), .ip2(n8618), .op(n5184) );
  nand3_1 U8778 ( .ip1(n8620), .ip2(miss), .ip3(cache_miss_count[0]), .op(
        n8621) );
  inv_1 U8779 ( .ip(cache_miss_count[1]), .op(n8622) );
  nor2_1 U8780 ( .ip1(n8621), .ip2(n8622), .op(n13228) );
  or2_1 U8781 ( .ip1(n8621), .ip2(n13228), .op(n8624) );
  or2_1 U8782 ( .ip1(n8622), .ip2(n13228), .op(n8623) );
  nand2_1 U8783 ( .ip1(n8624), .ip2(n8623), .op(n5190) );
  nand2_1 U8784 ( .ip1(n13228), .ip2(cache_miss_count[2]), .op(n13227) );
  inv_1 U8785 ( .ip(cache_miss_count[3]), .op(n8625) );
  nor2_1 U8786 ( .ip1(n13227), .ip2(n8625), .op(n13225) );
  or2_1 U8787 ( .ip1(n13227), .ip2(n13225), .op(n8627) );
  or2_1 U8788 ( .ip1(n8625), .ip2(n13225), .op(n8626) );
  nand2_1 U8789 ( .ip1(n8627), .ip2(n8626), .op(n5192) );
  inv_1 U8790 ( .ip(cache_miss_count[5]), .op(n8628) );
  nand2_1 U8791 ( .ip1(cache_miss_count[4]), .ip2(n13225), .op(n8629) );
  nor2_1 U8792 ( .ip1(n8628), .ip2(n8629), .op(n13222) );
  or2_1 U8793 ( .ip1(n8628), .ip2(n13222), .op(n8631) );
  or2_1 U8794 ( .ip1(n8629), .ip2(n13222), .op(n8630) );
  nand2_1 U8795 ( .ip1(n8631), .ip2(n8630), .op(n5194) );
  inv_1 U8796 ( .ip(cache_miss_count[8]), .op(n8632) );
  nand2_1 U8797 ( .ip1(n13222), .ip2(cache_miss_count[6]), .op(n13221) );
  inv_1 U8798 ( .ip(n13221), .op(n13224) );
  nand2_1 U8799 ( .ip1(n13224), .ip2(cache_miss_count[7]), .op(n8633) );
  nor2_1 U8800 ( .ip1(n8632), .ip2(n8633), .op(n13219) );
  or2_1 U8801 ( .ip1(n8632), .ip2(n13219), .op(n8635) );
  or2_1 U8802 ( .ip1(n8633), .ip2(n13219), .op(n8634) );
  nand2_1 U8803 ( .ip1(n8635), .ip2(n8634), .op(n5197) );
  inv_1 U8804 ( .ip(cache_miss_count[10]), .op(n8637) );
  nand4_1 U8805 ( .ip1(cache_miss_count[9]), .ip2(cache_miss_count[10]), .ip3(
        cache_miss_count[7]), .ip4(cache_miss_count[8]), .op(n8636) );
  nor2_1 U8806 ( .ip1(n13221), .ip2(n8636), .op(n13218) );
  or2_1 U8807 ( .ip1(n8637), .ip2(n13218), .op(n8640) );
  nand2_1 U8808 ( .ip1(cache_miss_count[9]), .ip2(n13219), .op(n8638) );
  or2_1 U8809 ( .ip1(n8638), .ip2(n13218), .op(n8639) );
  nand2_1 U8810 ( .ip1(n8640), .ip2(n8639), .op(n5199) );
  nand2_1 U8811 ( .ip1(n13218), .ip2(cache_miss_count[11]), .op(n8641) );
  inv_1 U8812 ( .ip(cache_miss_count[12]), .op(n8642) );
  nor2_1 U8813 ( .ip1(n8641), .ip2(n8642), .op(n13217) );
  or2_1 U8814 ( .ip1(n8641), .ip2(n13217), .op(n8644) );
  or2_1 U8815 ( .ip1(n8642), .ip2(n13217), .op(n8643) );
  nand2_1 U8816 ( .ip1(n8644), .ip2(n8643), .op(n5201) );
  nand2_1 U8817 ( .ip1(n13217), .ip2(cache_miss_count[13]), .op(n8645) );
  inv_1 U8818 ( .ip(cache_miss_count[14]), .op(n8646) );
  nor2_1 U8819 ( .ip1(n8645), .ip2(n8646), .op(n13216) );
  or2_1 U8820 ( .ip1(n8645), .ip2(n13216), .op(n8648) );
  or2_1 U8821 ( .ip1(n8646), .ip2(n13216), .op(n8647) );
  nand2_1 U8822 ( .ip1(n8648), .ip2(n8647), .op(n5203) );
  nand2_1 U8823 ( .ip1(n13216), .ip2(cache_miss_count[15]), .op(n8649) );
  inv_1 U8824 ( .ip(cache_miss_count[16]), .op(n8650) );
  nor2_1 U8825 ( .ip1(n8649), .ip2(n8650), .op(n13215) );
  or2_1 U8826 ( .ip1(n8649), .ip2(n13215), .op(n8652) );
  or2_1 U8827 ( .ip1(n8650), .ip2(n13215), .op(n8651) );
  nand2_1 U8828 ( .ip1(n8652), .ip2(n8651), .op(n5205) );
  nand2_1 U8829 ( .ip1(n13215), .ip2(cache_miss_count[17]), .op(n8653) );
  inv_1 U8830 ( .ip(cache_miss_count[18]), .op(n8654) );
  nor2_1 U8831 ( .ip1(n8653), .ip2(n8654), .op(n13214) );
  or2_1 U8832 ( .ip1(n8653), .ip2(n13214), .op(n8656) );
  or2_1 U8833 ( .ip1(n8654), .ip2(n13214), .op(n8655) );
  nand2_1 U8834 ( .ip1(n8656), .ip2(n8655), .op(n5207) );
  nand2_1 U8835 ( .ip1(n13214), .ip2(cache_miss_count[19]), .op(n8657) );
  inv_1 U8836 ( .ip(cache_miss_count[20]), .op(n8658) );
  nor2_1 U8837 ( .ip1(n8657), .ip2(n8658), .op(n13213) );
  or2_1 U8838 ( .ip1(n8657), .ip2(n13213), .op(n8660) );
  or2_1 U8839 ( .ip1(n8658), .ip2(n13213), .op(n8659) );
  nand2_1 U8840 ( .ip1(n8660), .ip2(n8659), .op(n5209) );
  nand2_1 U8841 ( .ip1(n13213), .ip2(cache_miss_count[21]), .op(n8661) );
  inv_1 U8842 ( .ip(cache_miss_count[22]), .op(n8662) );
  nor2_1 U8843 ( .ip1(n8661), .ip2(n8662), .op(n13212) );
  or2_1 U8844 ( .ip1(n8661), .ip2(n13212), .op(n8664) );
  or2_1 U8845 ( .ip1(n8662), .ip2(n13212), .op(n8663) );
  nand2_1 U8846 ( .ip1(n8664), .ip2(n8663), .op(n5211) );
  nand2_1 U8847 ( .ip1(n13212), .ip2(cache_miss_count[23]), .op(n8665) );
  inv_1 U8848 ( .ip(cache_miss_count[24]), .op(n8666) );
  nor2_1 U8849 ( .ip1(n8665), .ip2(n8666), .op(n13211) );
  or2_1 U8850 ( .ip1(n8665), .ip2(n13211), .op(n8668) );
  or2_1 U8851 ( .ip1(n8666), .ip2(n13211), .op(n8667) );
  nand2_1 U8852 ( .ip1(n8668), .ip2(n8667), .op(n5213) );
  nand2_1 U8853 ( .ip1(n13211), .ip2(cache_miss_count[25]), .op(n8669) );
  inv_1 U8854 ( .ip(cache_miss_count[26]), .op(n8670) );
  nor2_1 U8855 ( .ip1(n8669), .ip2(n8670), .op(n13210) );
  or2_1 U8856 ( .ip1(n8669), .ip2(n13210), .op(n8672) );
  or2_1 U8857 ( .ip1(n8670), .ip2(n13210), .op(n8671) );
  nand2_1 U8858 ( .ip1(n8672), .ip2(n8671), .op(n5215) );
  nand2_1 U8859 ( .ip1(n13210), .ip2(cache_miss_count[27]), .op(n8673) );
  inv_1 U8860 ( .ip(cache_miss_count[28]), .op(n8674) );
  nor2_1 U8861 ( .ip1(n8673), .ip2(n8674), .op(n13209) );
  or2_1 U8862 ( .ip1(n8673), .ip2(n13209), .op(n8676) );
  or2_1 U8863 ( .ip1(n8674), .ip2(n13209), .op(n8675) );
  nand2_1 U8864 ( .ip1(n8676), .ip2(n8675), .op(n5217) );
  inv_1 U8865 ( .ip(rst), .op(n13293) );
  buf_1 U8866 ( .ip(rst), .op(n12618) );
  inv_1 U8868 ( .ip(mem_data_cnt[3]), .op(n9701) );
  inv_1 U8869 ( .ip(mem_data_cnt[2]), .op(n9700) );
  nor2_1 U8870 ( .ip1(n9701), .ip2(n9700), .op(N4454) );
  inv_1 U8871 ( .ip(addr_req[8]), .op(n9162) );
  inv_1 U8872 ( .ip(addr_req[5]), .op(n8687) );
  inv_1 U8873 ( .ip(addr_req[6]), .op(n8679) );
  nand3_1 U8874 ( .ip1(n8687), .ip2(n8679), .ip3(addr_req[4]), .op(n8922) );
  inv_1 U8875 ( .ip(n8922), .op(n13278) );
  buf_1 U8876 ( .ip(n13278), .op(n9225) );
  nand2_1 U8877 ( .ip1(\cache_tag_A[1][1] ), .ip2(n9225), .op(n8690) );
  nor3_1 U8878 ( .ip1(addr_req[4]), .ip2(addr_req[5]), .ip3(addr_req[6]), .op(
        n13270) );
  nand3_1 U8879 ( .ip1(n8679), .ip2(addr_req[5]), .ip3(addr_req[4]), .op(
        n13266) );
  nor2_1 U8880 ( .ip1(n8677), .ip2(n13266), .op(n8686) );
  nand2_1 U8881 ( .ip1(addr_req[5]), .ip2(addr_req[6]), .op(n8678) );
  nor2_1 U8882 ( .ip1(addr_req[4]), .ip2(n8678), .op(n13251) );
  nand2_1 U8883 ( .ip1(\cache_tag_A[6][1] ), .ip2(n13251), .op(n8684) );
  nor3_1 U8884 ( .ip1(addr_req[4]), .ip2(addr_req[6]), .ip3(n8687), .op(n13264) );
  nand2_1 U8885 ( .ip1(\cache_tag_A[2][1] ), .ip2(n13264), .op(n8683) );
  inv_1 U8886 ( .ip(addr_req[4]), .op(n8680) );
  nand3_1 U8887 ( .ip1(n8680), .ip2(n8687), .ip3(addr_req[6]), .op(n8971) );
  inv_1 U8888 ( .ip(n8971), .op(n13268) );
  buf_1 U8889 ( .ip(n13268), .op(n9102) );
  nand2_1 U8890 ( .ip1(\cache_tag_A[4][1] ), .ip2(n9102), .op(n8682) );
  nor3_1 U8891 ( .ip1(n8680), .ip2(n8687), .ip3(n8679), .op(n13277) );
  nand2_1 U8892 ( .ip1(\cache_tag_A[7][1] ), .ip2(n13277), .op(n8681) );
  nand4_1 U8893 ( .ip1(n8684), .ip2(n8683), .ip3(n8682), .ip4(n8681), .op(
        n8685) );
  not_ab_or_c_or_d U8894 ( .ip1(n13270), .ip2(\cache_tag_A[0][1] ), .ip3(n8686), .ip4(n8685), .op(n8689) );
  nand3_1 U8895 ( .ip1(n8687), .ip2(addr_req[4]), .ip3(addr_req[6]), .op(n9164) );
  inv_1 U8896 ( .ip(n9164), .op(n13267) );
  nand2_1 U8897 ( .ip1(\cache_tag_A[5][1] ), .ip2(n13267), .op(n8688) );
  nand3_1 U8898 ( .ip1(n8690), .ip2(n8689), .ip3(n8688), .op(n8691) );
  mux2_1 U8899 ( .ip1(n9162), .ip2(addr_req[8]), .s(n8691), .op(n8730) );
  inv_1 U8900 ( .ip(addr_req[29]), .op(n9306) );
  nand2_1 U8901 ( .ip1(\cache_tag_A[6][22] ), .ip2(n13251), .op(n8701) );
  nor2_1 U8902 ( .ip1(n8692), .ip2(n9164), .op(n8698) );
  nand2_1 U8903 ( .ip1(\cache_tag_A[4][22] ), .ip2(n9102), .op(n8696) );
  nand2_1 U8904 ( .ip1(\cache_tag_A[7][22] ), .ip2(n13277), .op(n8695) );
  inv_1 U8905 ( .ip(n13266), .op(n13253) );
  buf_1 U8906 ( .ip(n13253), .op(n9271) );
  nand2_1 U8907 ( .ip1(\cache_tag_A[3][22] ), .ip2(n9271), .op(n8694) );
  nand2_1 U8908 ( .ip1(\cache_tag_A[1][22] ), .ip2(n9225), .op(n8693) );
  nand4_1 U8909 ( .ip1(n8696), .ip2(n8695), .ip3(n8694), .ip4(n8693), .op(
        n8697) );
  not_ab_or_c_or_d U8910 ( .ip1(n13270), .ip2(\cache_tag_A[0][22] ), .ip3(
        n8698), .ip4(n8697), .op(n8700) );
  nand2_1 U8911 ( .ip1(\cache_tag_A[2][22] ), .ip2(n13264), .op(n8699) );
  nand3_1 U8912 ( .ip1(n8701), .ip2(n8700), .ip3(n8699), .op(n8702) );
  mux2_1 U8913 ( .ip1(n9306), .ip2(addr_req[29]), .s(n8702), .op(n8729) );
  inv_1 U8914 ( .ip(addr_req[13]), .op(n8714) );
  nand2_1 U8915 ( .ip1(\cache_tag_A[5][6] ), .ip2(n13267), .op(n8712) );
  nor2_1 U8916 ( .ip1(n8703), .ip2(n8922), .op(n8709) );
  nand2_1 U8917 ( .ip1(\cache_tag_A[7][6] ), .ip2(n13277), .op(n8707) );
  nand2_1 U8918 ( .ip1(\cache_tag_A[2][6] ), .ip2(n13264), .op(n8706) );
  nand2_1 U8919 ( .ip1(\cache_tag_A[3][6] ), .ip2(n9271), .op(n8705) );
  nand2_1 U8920 ( .ip1(\cache_tag_A[0][6] ), .ip2(n13270), .op(n8704) );
  nand4_1 U8921 ( .ip1(n8707), .ip2(n8706), .ip3(n8705), .ip4(n8704), .op(
        n8708) );
  not_ab_or_c_or_d U8922 ( .ip1(n13251), .ip2(\cache_tag_A[6][6] ), .ip3(n8709), .ip4(n8708), .op(n8711) );
  nand2_1 U8923 ( .ip1(\cache_tag_A[4][6] ), .ip2(n9102), .op(n8710) );
  nand3_1 U8924 ( .ip1(n8712), .ip2(n8711), .ip3(n8710), .op(n8713) );
  mux2_1 U8925 ( .ip1(n8714), .ip2(addr_req[13]), .s(n8713), .op(n8728) );
  inv_1 U8926 ( .ip(addr_req[11]), .op(n8726) );
  nand2_1 U8927 ( .ip1(\cache_tag_A[1][4] ), .ip2(n9225), .op(n8724) );
  nor2_1 U8928 ( .ip1(n8715), .ip2(n13266), .op(n8721) );
  nand2_1 U8929 ( .ip1(\cache_tag_A[6][4] ), .ip2(n13251), .op(n8719) );
  nand2_1 U8930 ( .ip1(\cache_tag_A[0][4] ), .ip2(n13270), .op(n8718) );
  nand2_1 U8931 ( .ip1(\cache_tag_A[7][4] ), .ip2(n13277), .op(n8717) );
  nand2_1 U8932 ( .ip1(\cache_tag_A[5][4] ), .ip2(n13267), .op(n8716) );
  nand4_1 U8933 ( .ip1(n8719), .ip2(n8718), .ip3(n8717), .ip4(n8716), .op(
        n8720) );
  not_ab_or_c_or_d U8934 ( .ip1(n13268), .ip2(\cache_tag_A[4][4] ), .ip3(n8721), .ip4(n8720), .op(n8723) );
  nand2_1 U8935 ( .ip1(\cache_tag_A[2][4] ), .ip2(n13264), .op(n8722) );
  nand3_1 U8936 ( .ip1(n8724), .ip2(n8723), .ip3(n8722), .op(n8725) );
  mux2_1 U8937 ( .ip1(n8726), .ip2(addr_req[11]), .s(n8725), .op(n8727) );
  nand4_1 U8938 ( .ip1(n8730), .ip2(n8729), .ip3(n8728), .ip4(n8727), .op(
        n8994) );
  nand2_1 U8939 ( .ip1(\cache_tag_A[5][3] ), .ip2(n13267), .op(n8740) );
  buf_1 U8940 ( .ip(n13270), .op(n9165) );
  nor2_1 U8941 ( .ip1(n8731), .ip2(n8862), .op(n8737) );
  nand2_1 U8942 ( .ip1(\cache_tag_A[7][3] ), .ip2(n13277), .op(n8735) );
  nand2_1 U8943 ( .ip1(\cache_tag_A[4][3] ), .ip2(n9102), .op(n8734) );
  nand2_1 U8944 ( .ip1(\cache_tag_A[3][3] ), .ip2(n9271), .op(n8733) );
  nand2_1 U8945 ( .ip1(\cache_tag_A[1][3] ), .ip2(n9225), .op(n8732) );
  nand4_1 U8946 ( .ip1(n8735), .ip2(n8734), .ip3(n8733), .ip4(n8732), .op(
        n8736) );
  not_ab_or_c_or_d U8947 ( .ip1(n9165), .ip2(\cache_tag_A[0][3] ), .ip3(n8737), 
        .ip4(n8736), .op(n8739) );
  nand2_1 U8948 ( .ip1(\cache_tag_A[2][3] ), .ip2(n13264), .op(n8738) );
  nand3_1 U8949 ( .ip1(n8740), .ip2(n8739), .ip3(n8738), .op(n8741) );
  xor2_1 U8950 ( .ip1(addr_req[10]), .ip2(n8741), .op(n8993) );
  inv_1 U8951 ( .ip(addr_req[7]), .op(n8753) );
  nand2_1 U8952 ( .ip1(\cache_tag_A[3][0] ), .ip2(n9271), .op(n8751) );
  nand2_1 U8953 ( .ip1(\cache_tag_A[6][0] ), .ip2(n13251), .op(n8750) );
  nor2_1 U8954 ( .ip1(n8742), .ip2(n8922), .op(n8748) );
  nand2_1 U8955 ( .ip1(\cache_tag_A[2][0] ), .ip2(n13264), .op(n8746) );
  nand2_1 U8956 ( .ip1(\cache_tag_A[5][0] ), .ip2(n13267), .op(n8745) );
  nand2_1 U8957 ( .ip1(\cache_tag_A[0][0] ), .ip2(n13270), .op(n8744) );
  nand2_1 U8958 ( .ip1(\cache_tag_A[7][0] ), .ip2(n13277), .op(n8743) );
  nand4_1 U8959 ( .ip1(n8746), .ip2(n8745), .ip3(n8744), .ip4(n8743), .op(
        n8747) );
  not_ab_or_c_or_d U8960 ( .ip1(n13268), .ip2(\cache_tag_A[4][0] ), .ip3(n8748), .ip4(n8747), .op(n8749) );
  nand3_1 U8961 ( .ip1(n8751), .ip2(n8750), .ip3(n8749), .op(n8752) );
  mux2_1 U8962 ( .ip1(n8753), .ip2(addr_req[7]), .s(n8752), .op(n8791) );
  inv_1 U8963 ( .ip(addr_req[19]), .op(n9189) );
  nand2_1 U8964 ( .ip1(\cache_tag_A[2][12] ), .ip2(n13264), .op(n8763) );
  nor2_1 U8965 ( .ip1(n8754), .ip2(n8971), .op(n8760) );
  nand2_1 U8966 ( .ip1(\cache_tag_A[3][12] ), .ip2(n9271), .op(n8758) );
  nand2_1 U8967 ( .ip1(\cache_tag_A[7][12] ), .ip2(n13277), .op(n8757) );
  nand2_1 U8968 ( .ip1(\cache_tag_A[1][12] ), .ip2(n9225), .op(n8756) );
  nand2_1 U8969 ( .ip1(\cache_tag_A[5][12] ), .ip2(n13267), .op(n8755) );
  nand4_1 U8970 ( .ip1(n8758), .ip2(n8757), .ip3(n8756), .ip4(n8755), .op(
        n8759) );
  not_ab_or_c_or_d U8971 ( .ip1(n13251), .ip2(\cache_tag_A[6][12] ), .ip3(
        n8760), .ip4(n8759), .op(n8762) );
  nand2_1 U8972 ( .ip1(\cache_tag_A[0][12] ), .ip2(n9165), .op(n8761) );
  nand3_1 U8973 ( .ip1(n8763), .ip2(n8762), .ip3(n8761), .op(n8764) );
  mux2_1 U8974 ( .ip1(n9189), .ip2(addr_req[19]), .s(n8764), .op(n8790) );
  inv_1 U8975 ( .ip(addr_req[12]), .op(n8776) );
  nand2_1 U8976 ( .ip1(\cache_tag_A[1][5] ), .ip2(n9225), .op(n8774) );
  nor2_1 U8977 ( .ip1(n8765), .ip2(n9164), .op(n8771) );
  nand2_1 U8978 ( .ip1(\cache_tag_A[7][5] ), .ip2(n13277), .op(n8769) );
  nand2_1 U8979 ( .ip1(\cache_tag_A[6][5] ), .ip2(n13251), .op(n8768) );
  nand2_1 U8980 ( .ip1(\cache_tag_A[2][5] ), .ip2(n13264), .op(n8767) );
  nand2_1 U8981 ( .ip1(\cache_tag_A[4][5] ), .ip2(n9102), .op(n8766) );
  nand4_1 U8982 ( .ip1(n8769), .ip2(n8768), .ip3(n8767), .ip4(n8766), .op(
        n8770) );
  not_ab_or_c_or_d U8983 ( .ip1(n13253), .ip2(\cache_tag_A[3][5] ), .ip3(n8771), .ip4(n8770), .op(n8773) );
  nand2_1 U8984 ( .ip1(\cache_tag_A[0][5] ), .ip2(n9165), .op(n8772) );
  nand3_1 U8985 ( .ip1(n8774), .ip2(n8773), .ip3(n8772), .op(n8775) );
  mux2_1 U8986 ( .ip1(n8776), .ip2(addr_req[12]), .s(n8775), .op(n8789) );
  inv_1 U8987 ( .ip(addr_req[22]), .op(n9217) );
  nand2_1 U8988 ( .ip1(\cache_tag_A[0][15] ), .ip2(n9165), .op(n8786) );
  nor2_1 U8989 ( .ip1(n8777), .ip2(n13266), .op(n8783) );
  nand2_1 U8990 ( .ip1(\cache_tag_A[6][15] ), .ip2(n13251), .op(n8781) );
  nand2_1 U8991 ( .ip1(\cache_tag_A[7][15] ), .ip2(n13277), .op(n8780) );
  nand2_1 U8992 ( .ip1(\cache_tag_A[1][15] ), .ip2(n9225), .op(n8779) );
  nand2_1 U8993 ( .ip1(\cache_tag_A[4][15] ), .ip2(n9102), .op(n8778) );
  nand4_1 U8994 ( .ip1(n8781), .ip2(n8780), .ip3(n8779), .ip4(n8778), .op(
        n8782) );
  not_ab_or_c_or_d U8995 ( .ip1(n13264), .ip2(\cache_tag_A[2][15] ), .ip3(
        n8783), .ip4(n8782), .op(n8785) );
  nand2_1 U8996 ( .ip1(\cache_tag_A[5][15] ), .ip2(n13267), .op(n8784) );
  nand3_1 U8997 ( .ip1(n8786), .ip2(n8785), .ip3(n8784), .op(n8787) );
  mux2_1 U8998 ( .ip1(n9217), .ip2(addr_req[22]), .s(n8787), .op(n8788) );
  nand4_1 U8999 ( .ip1(n8791), .ip2(n8790), .ip3(n8789), .ip4(n8788), .op(
        n8992) );
  nand2_1 U9000 ( .ip1(\cache_tag_A[0][11] ), .ip2(n13270), .op(n8801) );
  nor2_1 U9001 ( .ip1(n8792), .ip2(n8862), .op(n8798) );
  nand2_1 U9002 ( .ip1(\cache_tag_A[7][11] ), .ip2(n13277), .op(n8796) );
  nand2_1 U9003 ( .ip1(\cache_tag_A[4][11] ), .ip2(n9102), .op(n8795) );
  buf_1 U9004 ( .ip(n13264), .op(n9349) );
  nand2_1 U9005 ( .ip1(\cache_tag_A[2][11] ), .ip2(n9349), .op(n8794) );
  nand2_1 U9006 ( .ip1(\cache_tag_A[3][11] ), .ip2(n9271), .op(n8793) );
  nand4_1 U9007 ( .ip1(n8796), .ip2(n8795), .ip3(n8794), .ip4(n8793), .op(
        n8797) );
  not_ab_or_c_or_d U9008 ( .ip1(n13278), .ip2(\cache_tag_A[1][11] ), .ip3(
        n8798), .ip4(n8797), .op(n8800) );
  nand2_1 U9009 ( .ip1(\cache_tag_A[5][11] ), .ip2(n13267), .op(n8799) );
  nand3_1 U9010 ( .ip1(n8801), .ip2(n8800), .ip3(n8799), .op(n8802) );
  xor2_1 U9011 ( .ip1(addr_req[18]), .ip2(n8802), .op(n8839) );
  nand2_1 U9012 ( .ip1(\cache_tag_A[5][10] ), .ip2(n13267), .op(n8812) );
  nand2_1 U9013 ( .ip1(\cache_tag_A[2][10] ), .ip2(n13264), .op(n8811) );
  nor2_1 U9014 ( .ip1(n8803), .ip2(n13266), .op(n8809) );
  nand2_1 U9015 ( .ip1(\cache_tag_A[6][10] ), .ip2(n13251), .op(n8807) );
  nand2_1 U9016 ( .ip1(\cache_tag_A[1][10] ), .ip2(n9225), .op(n8806) );
  nand2_1 U9017 ( .ip1(\cache_tag_A[0][10] ), .ip2(n13270), .op(n8805) );
  nand2_1 U9018 ( .ip1(\cache_tag_A[7][10] ), .ip2(n13277), .op(n8804) );
  nand4_1 U9019 ( .ip1(n8807), .ip2(n8806), .ip3(n8805), .ip4(n8804), .op(
        n8808) );
  not_ab_or_c_or_d U9020 ( .ip1(n9102), .ip2(\cache_tag_A[4][10] ), .ip3(n8809), .ip4(n8808), .op(n8810) );
  nand3_1 U9021 ( .ip1(n8812), .ip2(n8811), .ip3(n8810), .op(n8813) );
  xor2_1 U9022 ( .ip1(addr_req[17]), .ip2(n8813), .op(n8838) );
  nand2_1 U9023 ( .ip1(\cache_tag_A[7][9] ), .ip2(n13277), .op(n8823) );
  buf_1 U9024 ( .ip(n13267), .op(n13254) );
  nor2_1 U9025 ( .ip1(n8814), .ip2(n8971), .op(n8820) );
  nand2_1 U9026 ( .ip1(\cache_tag_A[3][9] ), .ip2(n9271), .op(n8818) );
  nand2_1 U9027 ( .ip1(\cache_tag_A[6][9] ), .ip2(n13251), .op(n8817) );
  nand2_1 U9028 ( .ip1(\cache_tag_A[1][9] ), .ip2(n9225), .op(n8816) );
  nand2_1 U9029 ( .ip1(\cache_tag_A[0][9] ), .ip2(n13270), .op(n8815) );
  nand4_1 U9030 ( .ip1(n8818), .ip2(n8817), .ip3(n8816), .ip4(n8815), .op(
        n8819) );
  not_ab_or_c_or_d U9031 ( .ip1(n13254), .ip2(\cache_tag_A[5][9] ), .ip3(n8820), .ip4(n8819), .op(n8822) );
  nand2_1 U9032 ( .ip1(\cache_tag_A[2][9] ), .ip2(n13264), .op(n8821) );
  nand3_1 U9033 ( .ip1(n8823), .ip2(n8822), .ip3(n8821), .op(n8824) );
  xor2_1 U9034 ( .ip1(addr_req[16]), .ip2(n8824), .op(n8837) );
  nand2_1 U9035 ( .ip1(\cache_tag_A[7][8] ), .ip2(n13277), .op(n8834) );
  inv_1 U9036 ( .ip(n13251), .op(n8862) );
  nor2_1 U9037 ( .ip1(n8825), .ip2(n8862), .op(n8831) );
  nand2_1 U9038 ( .ip1(\cache_tag_A[4][8] ), .ip2(n9102), .op(n8829) );
  nand2_1 U9039 ( .ip1(\cache_tag_A[2][8] ), .ip2(n9349), .op(n8828) );
  nand2_1 U9040 ( .ip1(\cache_tag_A[3][8] ), .ip2(n9271), .op(n8827) );
  nand2_1 U9041 ( .ip1(\cache_tag_A[0][8] ), .ip2(n13270), .op(n8826) );
  nand4_1 U9042 ( .ip1(n8829), .ip2(n8828), .ip3(n8827), .ip4(n8826), .op(
        n8830) );
  not_ab_or_c_or_d U9043 ( .ip1(n13254), .ip2(\cache_tag_A[5][8] ), .ip3(n8831), .ip4(n8830), .op(n8833) );
  nand2_1 U9044 ( .ip1(\cache_tag_A[1][8] ), .ip2(n9225), .op(n8832) );
  nand3_1 U9045 ( .ip1(n8834), .ip2(n8833), .ip3(n8832), .op(n8835) );
  xor2_1 U9046 ( .ip1(addr_req[15]), .ip2(n8835), .op(n8836) );
  nor4_1 U9047 ( .ip1(n8839), .ip2(n8838), .ip3(n8837), .ip4(n8836), .op(n8990) );
  nand2_1 U9048 ( .ip1(\cache_tag_A[3][18] ), .ip2(n9271), .op(n8849) );
  nor2_1 U9049 ( .ip1(n8840), .ip2(n8971), .op(n8846) );
  nand2_1 U9050 ( .ip1(\cache_tag_A[7][18] ), .ip2(n13277), .op(n8844) );
  nand2_1 U9051 ( .ip1(\cache_tag_A[2][18] ), .ip2(n13264), .op(n8843) );
  nand2_1 U9052 ( .ip1(\cache_tag_A[5][18] ), .ip2(n13267), .op(n8842) );
  nand2_1 U9053 ( .ip1(\cache_tag_A[0][18] ), .ip2(n13270), .op(n8841) );
  nand4_1 U9054 ( .ip1(n8844), .ip2(n8843), .ip3(n8842), .ip4(n8841), .op(
        n8845) );
  not_ab_or_c_or_d U9055 ( .ip1(n13278), .ip2(\cache_tag_A[1][18] ), .ip3(
        n8846), .ip4(n8845), .op(n8848) );
  nand2_1 U9056 ( .ip1(\cache_tag_A[6][18] ), .ip2(n13251), .op(n8847) );
  nand3_1 U9057 ( .ip1(n8849), .ip2(n8848), .ip3(n8847), .op(n8850) );
  xor2_1 U9058 ( .ip1(addr_req[25]), .ip2(n8850), .op(n8888) );
  nand2_1 U9059 ( .ip1(\cache_tag_A[2][7] ), .ip2(n13264), .op(n8860) );
  nor2_1 U9060 ( .ip1(n8851), .ip2(n8971), .op(n8857) );
  nand2_1 U9061 ( .ip1(\cache_tag_A[5][7] ), .ip2(n13267), .op(n8855) );
  nand2_1 U9062 ( .ip1(\cache_tag_A[3][7] ), .ip2(n9271), .op(n8854) );
  nand2_1 U9063 ( .ip1(\cache_tag_A[1][7] ), .ip2(n9225), .op(n8853) );
  nand2_1 U9064 ( .ip1(\cache_tag_A[7][7] ), .ip2(n13277), .op(n8852) );
  nand4_1 U9065 ( .ip1(n8855), .ip2(n8854), .ip3(n8853), .ip4(n8852), .op(
        n8856) );
  not_ab_or_c_or_d U9066 ( .ip1(n9165), .ip2(\cache_tag_A[0][7] ), .ip3(n8857), 
        .ip4(n8856), .op(n8859) );
  nand2_1 U9067 ( .ip1(\cache_tag_A[6][7] ), .ip2(n13251), .op(n8858) );
  nand3_1 U9068 ( .ip1(n8860), .ip2(n8859), .ip3(n8858), .op(n8861) );
  xor2_1 U9069 ( .ip1(addr_req[14]), .ip2(n8861), .op(n8887) );
  nand2_1 U9070 ( .ip1(\cache_tag_A[2][21] ), .ip2(n13264), .op(n8872) );
  nor2_1 U9071 ( .ip1(n8863), .ip2(n8862), .op(n8869) );
  nand2_1 U9072 ( .ip1(\cache_tag_A[3][21] ), .ip2(n9271), .op(n8867) );
  nand2_1 U9073 ( .ip1(\cache_tag_A[0][21] ), .ip2(n9165), .op(n8866) );
  nand2_1 U9074 ( .ip1(\cache_tag_A[1][21] ), .ip2(n9225), .op(n8865) );
  nand2_1 U9075 ( .ip1(\cache_tag_A[7][21] ), .ip2(n13277), .op(n8864) );
  nand4_1 U9076 ( .ip1(n8867), .ip2(n8866), .ip3(n8865), .ip4(n8864), .op(
        n8868) );
  not_ab_or_c_or_d U9077 ( .ip1(n9102), .ip2(\cache_tag_A[4][21] ), .ip3(n8869), .ip4(n8868), .op(n8871) );
  nand2_1 U9078 ( .ip1(\cache_tag_A[5][21] ), .ip2(n13267), .op(n8870) );
  nand3_1 U9079 ( .ip1(n8872), .ip2(n8871), .ip3(n8870), .op(n8873) );
  xor2_1 U9080 ( .ip1(addr_req[28]), .ip2(n8873), .op(n8886) );
  nand2_1 U9081 ( .ip1(\cache_tag_A[2][16] ), .ip2(n13264), .op(n8883) );
  nor2_1 U9082 ( .ip1(n8874), .ip2(n9164), .op(n8880) );
  nand2_1 U9083 ( .ip1(\cache_tag_A[1][16] ), .ip2(n13278), .op(n8878) );
  nand2_1 U9084 ( .ip1(\cache_tag_A[4][16] ), .ip2(n9102), .op(n8877) );
  nand2_1 U9085 ( .ip1(\cache_tag_A[6][16] ), .ip2(n13251), .op(n8876) );
  nand2_1 U9086 ( .ip1(\cache_tag_A[3][16] ), .ip2(n9271), .op(n8875) );
  nand4_1 U9087 ( .ip1(n8878), .ip2(n8877), .ip3(n8876), .ip4(n8875), .op(
        n8879) );
  not_ab_or_c_or_d U9088 ( .ip1(n13277), .ip2(\cache_tag_A[7][16] ), .ip3(
        n8880), .ip4(n8879), .op(n8882) );
  nand2_1 U9089 ( .ip1(\cache_tag_A[0][16] ), .ip2(n13270), .op(n8881) );
  nand3_1 U9090 ( .ip1(n8883), .ip2(n8882), .ip3(n8881), .op(n8884) );
  xor2_1 U9091 ( .ip1(addr_req[23]), .ip2(n8884), .op(n8885) );
  nor4_1 U9092 ( .ip1(n8888), .ip2(n8887), .ip3(n8886), .ip4(n8885), .op(n8989) );
  nand2_1 U9093 ( .ip1(\cache_tag_A[1][17] ), .ip2(n13278), .op(n8898) );
  buf_1 U9094 ( .ip(n13251), .op(n13269) );
  nor2_1 U9095 ( .ip1(n8889), .ip2(n8971), .op(n8895) );
  nand2_1 U9096 ( .ip1(\cache_tag_A[3][17] ), .ip2(n9271), .op(n8893) );
  nand2_1 U9097 ( .ip1(\cache_tag_A[7][17] ), .ip2(n13277), .op(n8892) );
  nand2_1 U9098 ( .ip1(\cache_tag_A[5][17] ), .ip2(n13254), .op(n8891) );
  nand2_1 U9099 ( .ip1(\cache_tag_A[2][17] ), .ip2(n13264), .op(n8890) );
  nand4_1 U9100 ( .ip1(n8893), .ip2(n8892), .ip3(n8891), .ip4(n8890), .op(
        n8894) );
  not_ab_or_c_or_d U9101 ( .ip1(n13269), .ip2(\cache_tag_A[6][17] ), .ip3(
        n8895), .ip4(n8894), .op(n8897) );
  nand2_1 U9102 ( .ip1(\cache_tag_A[0][17] ), .ip2(n13270), .op(n8896) );
  nand3_1 U9103 ( .ip1(n8898), .ip2(n8897), .ip3(n8896), .op(n8899) );
  xor2_1 U9104 ( .ip1(addr_req[24]), .ip2(n8899), .op(n8937) );
  nand2_1 U9105 ( .ip1(\cache_tag_A[2][24] ), .ip2(n13264), .op(n8909) );
  nor2_1 U9106 ( .ip1(n8900), .ip2(n8922), .op(n8906) );
  nand2_1 U9107 ( .ip1(\cache_tag_A[5][24] ), .ip2(n13254), .op(n8904) );
  nand2_1 U9108 ( .ip1(\cache_tag_A[7][24] ), .ip2(n13277), .op(n8903) );
  nand2_1 U9109 ( .ip1(\cache_tag_A[3][24] ), .ip2(n13253), .op(n8902) );
  nand2_1 U9110 ( .ip1(\cache_tag_A[6][24] ), .ip2(n13251), .op(n8901) );
  nand4_1 U9111 ( .ip1(n8904), .ip2(n8903), .ip3(n8902), .ip4(n8901), .op(
        n8905) );
  not_ab_or_c_or_d U9112 ( .ip1(n9102), .ip2(\cache_tag_A[4][24] ), .ip3(n8906), .ip4(n8905), .op(n8908) );
  nand2_1 U9113 ( .ip1(\cache_tag_A[0][24] ), .ip2(n13270), .op(n8907) );
  nand3_1 U9114 ( .ip1(n8909), .ip2(n8908), .ip3(n8907), .op(n8910) );
  xor2_1 U9115 ( .ip1(addr_req[31]), .ip2(n8910), .op(n8936) );
  nand2_1 U9116 ( .ip1(\cache_tag_A[2][13] ), .ip2(n13264), .op(n8920) );
  nor2_1 U9117 ( .ip1(n8911), .ip2(n9164), .op(n8917) );
  nand2_1 U9118 ( .ip1(\cache_tag_A[4][13] ), .ip2(n9102), .op(n8915) );
  nand2_1 U9119 ( .ip1(\cache_tag_A[0][13] ), .ip2(n9165), .op(n8914) );
  nand2_1 U9120 ( .ip1(\cache_tag_A[6][13] ), .ip2(n13251), .op(n8913) );
  nand2_1 U9121 ( .ip1(\cache_tag_A[7][13] ), .ip2(n13277), .op(n8912) );
  nand4_1 U9122 ( .ip1(n8915), .ip2(n8914), .ip3(n8913), .ip4(n8912), .op(
        n8916) );
  not_ab_or_c_or_d U9123 ( .ip1(n13278), .ip2(\cache_tag_A[1][13] ), .ip3(
        n8917), .ip4(n8916), .op(n8919) );
  nand2_1 U9124 ( .ip1(\cache_tag_A[3][13] ), .ip2(n13253), .op(n8918) );
  nand3_1 U9125 ( .ip1(n8920), .ip2(n8919), .ip3(n8918), .op(n8921) );
  xor2_1 U9126 ( .ip1(addr_req[20]), .ip2(n8921), .op(n8935) );
  nand2_1 U9127 ( .ip1(\cache_tag_A[6][19] ), .ip2(n13251), .op(n8932) );
  nor2_1 U9128 ( .ip1(n8923), .ip2(n8922), .op(n8929) );
  nand2_1 U9129 ( .ip1(\cache_tag_A[4][19] ), .ip2(n9102), .op(n8927) );
  nand2_1 U9130 ( .ip1(\cache_tag_A[2][19] ), .ip2(n9349), .op(n8926) );
  nand2_1 U9131 ( .ip1(\cache_tag_A[5][19] ), .ip2(n13254), .op(n8925) );
  nand2_1 U9132 ( .ip1(\cache_tag_A[3][19] ), .ip2(n9271), .op(n8924) );
  nand4_1 U9133 ( .ip1(n8927), .ip2(n8926), .ip3(n8925), .ip4(n8924), .op(
        n8928) );
  not_ab_or_c_or_d U9134 ( .ip1(n13277), .ip2(\cache_tag_A[7][19] ), .ip3(
        n8929), .ip4(n8928), .op(n8931) );
  nand2_1 U9135 ( .ip1(\cache_tag_A[0][19] ), .ip2(n13270), .op(n8930) );
  nand3_1 U9136 ( .ip1(n8932), .ip2(n8931), .ip3(n8930), .op(n8933) );
  xor2_1 U9137 ( .ip1(addr_req[26]), .ip2(n8933), .op(n8934) );
  nor4_1 U9138 ( .ip1(n8937), .ip2(n8936), .ip3(n8935), .ip4(n8934), .op(n8988) );
  nand2_1 U9139 ( .ip1(\cache_tag_A[7][14] ), .ip2(n13277), .op(n8947) );
  nor2_1 U9140 ( .ip1(n8938), .ip2(n13266), .op(n8944) );
  nand2_1 U9141 ( .ip1(\cache_tag_A[1][14] ), .ip2(n13278), .op(n8942) );
  nand2_1 U9142 ( .ip1(\cache_tag_A[2][14] ), .ip2(n13264), .op(n8941) );
  nand2_1 U9143 ( .ip1(\cache_tag_A[4][14] ), .ip2(n13268), .op(n8940) );
  nand2_1 U9144 ( .ip1(\cache_tag_A[0][14] ), .ip2(n13270), .op(n8939) );
  nand4_1 U9145 ( .ip1(n8942), .ip2(n8941), .ip3(n8940), .ip4(n8939), .op(
        n8943) );
  not_ab_or_c_or_d U9146 ( .ip1(n13269), .ip2(\cache_tag_A[6][14] ), .ip3(
        n8944), .ip4(n8943), .op(n8946) );
  nand2_1 U9147 ( .ip1(\cache_tag_A[5][14] ), .ip2(n13254), .op(n8945) );
  nand3_1 U9148 ( .ip1(n8947), .ip2(n8946), .ip3(n8945), .op(n8948) );
  xor2_1 U9149 ( .ip1(addr_req[21]), .ip2(n8948), .op(n8986) );
  nand2_1 U9150 ( .ip1(\cache_tag_A[4][23] ), .ip2(n9102), .op(n8958) );
  nor2_1 U9151 ( .ip1(n8949), .ip2(n9178), .op(n8955) );
  nand2_1 U9152 ( .ip1(\cache_tag_A[5][23] ), .ip2(n13254), .op(n8953) );
  nand2_1 U9153 ( .ip1(\cache_tag_A[3][23] ), .ip2(n13253), .op(n8952) );
  nand2_1 U9154 ( .ip1(\cache_tag_A[1][23] ), .ip2(n9225), .op(n8951) );
  nand2_1 U9155 ( .ip1(\cache_tag_A[2][23] ), .ip2(n13264), .op(n8950) );
  nand4_1 U9156 ( .ip1(n8953), .ip2(n8952), .ip3(n8951), .ip4(n8950), .op(
        n8954) );
  not_ab_or_c_or_d U9157 ( .ip1(n9165), .ip2(\cache_tag_A[0][23] ), .ip3(n8955), .ip4(n8954), .op(n8957) );
  nand2_1 U9158 ( .ip1(\cache_tag_A[6][23] ), .ip2(n13251), .op(n8956) );
  nand3_1 U9159 ( .ip1(n8958), .ip2(n8957), .ip3(n8956), .op(n8959) );
  xor2_1 U9160 ( .ip1(addr_req[30]), .ip2(n8959), .op(n8985) );
  nand2_1 U9161 ( .ip1(\cache_tag_A[0][2] ), .ip2(n13270), .op(n8969) );
  nor2_1 U9162 ( .ip1(n8960), .ip2(n9164), .op(n8966) );
  nand2_1 U9163 ( .ip1(\cache_tag_A[6][2] ), .ip2(n13251), .op(n8964) );
  nand2_1 U9164 ( .ip1(\cache_tag_A[7][2] ), .ip2(n13277), .op(n8963) );
  nand2_1 U9165 ( .ip1(\cache_tag_A[4][2] ), .ip2(n9102), .op(n8962) );
  nand2_1 U9166 ( .ip1(\cache_tag_A[3][2] ), .ip2(n13253), .op(n8961) );
  nand4_1 U9167 ( .ip1(n8964), .ip2(n8963), .ip3(n8962), .ip4(n8961), .op(
        n8965) );
  not_ab_or_c_or_d U9168 ( .ip1(n9349), .ip2(\cache_tag_A[2][2] ), .ip3(n8966), 
        .ip4(n8965), .op(n8968) );
  nand2_1 U9169 ( .ip1(\cache_tag_A[1][2] ), .ip2(n9225), .op(n8967) );
  nand3_1 U9170 ( .ip1(n8969), .ip2(n8968), .ip3(n8967), .op(n8970) );
  xor2_1 U9171 ( .ip1(addr_req[9]), .ip2(n8970), .op(n8984) );
  nand2_1 U9172 ( .ip1(\cache_tag_A[0][20] ), .ip2(n13270), .op(n8981) );
  nor2_1 U9173 ( .ip1(n8972), .ip2(n8971), .op(n8978) );
  nand2_1 U9174 ( .ip1(\cache_tag_A[1][20] ), .ip2(n13278), .op(n8976) );
  nand2_1 U9175 ( .ip1(\cache_tag_A[3][20] ), .ip2(n13253), .op(n8975) );
  nand2_1 U9176 ( .ip1(\cache_tag_A[6][20] ), .ip2(n13251), .op(n8974) );
  nand2_1 U9177 ( .ip1(\cache_tag_A[7][20] ), .ip2(n13277), .op(n8973) );
  nand4_1 U9178 ( .ip1(n8976), .ip2(n8975), .ip3(n8974), .ip4(n8973), .op(
        n8977) );
  not_ab_or_c_or_d U9179 ( .ip1(n13254), .ip2(\cache_tag_A[5][20] ), .ip3(
        n8978), .ip4(n8977), .op(n8980) );
  nand2_1 U9180 ( .ip1(\cache_tag_A[2][20] ), .ip2(n13264), .op(n8979) );
  nand3_1 U9181 ( .ip1(n8981), .ip2(n8980), .ip3(n8979), .op(n8982) );
  xor2_1 U9182 ( .ip1(addr_req[27]), .ip2(n8982), .op(n8983) );
  nor4_1 U9183 ( .ip1(n8986), .ip2(n8985), .ip3(n8984), .ip4(n8983), .op(n8987) );
  nand4_1 U9184 ( .ip1(n8990), .ip2(n8989), .ip3(n8988), .ip4(n8987), .op(
        n8991) );
  nor4_1 U9185 ( .ip1(n8994), .ip2(n8993), .ip3(n8992), .ip4(n8991), .op(
        n13283) );
  nand2_1 U9186 ( .ip1(\cache_tag_B[3][3] ), .ip2(n13253), .op(n9004) );
  nor2_1 U9187 ( .ip1(n9178), .ip2(n8995), .op(n9001) );
  nand2_1 U9188 ( .ip1(n13267), .ip2(\cache_tag_B[5][3] ), .op(n8999) );
  nand2_1 U9189 ( .ip1(n13268), .ip2(\cache_tag_B[4][3] ), .op(n8998) );
  nand2_1 U9190 ( .ip1(n9165), .ip2(\cache_tag_B[0][3] ), .op(n8997) );
  nand2_1 U9191 ( .ip1(n13264), .ip2(\cache_tag_B[2][3] ), .op(n8996) );
  nand4_1 U9192 ( .ip1(n8999), .ip2(n8998), .ip3(n8997), .ip4(n8996), .op(
        n9000) );
  not_ab_or_c_or_d U9193 ( .ip1(n13251), .ip2(\cache_tag_B[6][3] ), .ip3(n9001), .ip4(n9000), .op(n9003) );
  nand2_1 U9194 ( .ip1(n13278), .ip2(\cache_tag_B[1][3] ), .op(n9002) );
  nand3_1 U9195 ( .ip1(n9004), .ip2(n9003), .ip3(n9002), .op(n9005) );
  xor2_1 U9196 ( .ip1(addr_req[10]), .ip2(n9005), .op(n9042) );
  nand2_1 U9197 ( .ip1(\cache_tag_B[2][20] ), .ip2(n13264), .op(n9015) );
  nor2_1 U9198 ( .ip1(n9178), .ip2(n9006), .op(n9012) );
  nand2_1 U9199 ( .ip1(n13270), .ip2(\cache_tag_B[0][20] ), .op(n9010) );
  nand2_1 U9200 ( .ip1(n13268), .ip2(\cache_tag_B[4][20] ), .op(n9009) );
  nand2_1 U9201 ( .ip1(n13253), .ip2(\cache_tag_B[3][20] ), .op(n9008) );
  nand2_1 U9202 ( .ip1(n13267), .ip2(\cache_tag_B[5][20] ), .op(n9007) );
  nand4_1 U9203 ( .ip1(n9010), .ip2(n9009), .ip3(n9008), .ip4(n9007), .op(
        n9011) );
  not_ab_or_c_or_d U9204 ( .ip1(n13251), .ip2(\cache_tag_B[6][20] ), .ip3(
        n9012), .ip4(n9011), .op(n9014) );
  nand2_1 U9205 ( .ip1(n13278), .ip2(\cache_tag_B[1][20] ), .op(n9013) );
  nand3_1 U9206 ( .ip1(n9015), .ip2(n9014), .ip3(n9013), .op(n9016) );
  xor2_1 U9207 ( .ip1(addr_req[27]), .ip2(n9016), .op(n9041) );
  nand2_1 U9208 ( .ip1(n13251), .ip2(\cache_tag_B[6][5] ), .op(n9026) );
  nor2_1 U9209 ( .ip1(n9164), .ip2(n9017), .op(n9023) );
  nand2_1 U9210 ( .ip1(n13270), .ip2(\cache_tag_B[0][5] ), .op(n9021) );
  nand2_1 U9211 ( .ip1(n13278), .ip2(\cache_tag_B[1][5] ), .op(n9020) );
  nand2_1 U9212 ( .ip1(n13277), .ip2(\cache_tag_B[7][5] ), .op(n9019) );
  nand2_1 U9213 ( .ip1(n13268), .ip2(\cache_tag_B[4][5] ), .op(n9018) );
  nand4_1 U9214 ( .ip1(n9021), .ip2(n9020), .ip3(n9019), .ip4(n9018), .op(
        n9022) );
  not_ab_or_c_or_d U9215 ( .ip1(\cache_tag_B[3][5] ), .ip2(n13253), .ip3(n9023), .ip4(n9022), .op(n9025) );
  nand2_1 U9216 ( .ip1(n13264), .ip2(\cache_tag_B[2][5] ), .op(n9024) );
  nand3_1 U9217 ( .ip1(n9026), .ip2(n9025), .ip3(n9024), .op(n9027) );
  xor2_1 U9218 ( .ip1(addr_req[12]), .ip2(n9027), .op(n9040) );
  nand2_1 U9219 ( .ip1(\cache_tag_B[6][18] ), .ip2(n13251), .op(n9037) );
  nor2_1 U9220 ( .ip1(n9178), .ip2(n9028), .op(n9034) );
  nand2_1 U9221 ( .ip1(n13268), .ip2(\cache_tag_B[4][18] ), .op(n9032) );
  nand2_1 U9222 ( .ip1(n13270), .ip2(\cache_tag_B[0][18] ), .op(n9031) );
  nand2_1 U9223 ( .ip1(n13264), .ip2(\cache_tag_B[2][18] ), .op(n9030) );
  nand2_1 U9224 ( .ip1(n13253), .ip2(\cache_tag_B[3][18] ), .op(n9029) );
  nand4_1 U9225 ( .ip1(n9032), .ip2(n9031), .ip3(n9030), .ip4(n9029), .op(
        n9033) );
  not_ab_or_c_or_d U9226 ( .ip1(n13254), .ip2(\cache_tag_B[5][18] ), .ip3(
        n9034), .ip4(n9033), .op(n9036) );
  nand2_1 U9227 ( .ip1(n13278), .ip2(\cache_tag_B[1][18] ), .op(n9035) );
  nand3_1 U9228 ( .ip1(n9037), .ip2(n9036), .ip3(n9035), .op(n9038) );
  xor2_1 U9229 ( .ip1(addr_req[25]), .ip2(n9038), .op(n9039) );
  nor4_1 U9230 ( .ip1(n9042), .ip2(n9041), .ip3(n9040), .ip4(n9039), .op(n9318) );
  nand2_1 U9231 ( .ip1(\cache_tag_B[2][6] ), .ip2(n13264), .op(n9052) );
  nor2_1 U9232 ( .ip1(n9178), .ip2(n9043), .op(n9049) );
  nand2_1 U9233 ( .ip1(n13269), .ip2(\cache_tag_B[6][6] ), .op(n9047) );
  nand2_1 U9234 ( .ip1(n13254), .ip2(\cache_tag_B[5][6] ), .op(n9046) );
  nand2_1 U9235 ( .ip1(n13270), .ip2(\cache_tag_B[0][6] ), .op(n9045) );
  nand2_1 U9236 ( .ip1(n13268), .ip2(\cache_tag_B[4][6] ), .op(n9044) );
  nand4_1 U9237 ( .ip1(n9047), .ip2(n9046), .ip3(n9045), .ip4(n9044), .op(
        n9048) );
  not_ab_or_c_or_d U9238 ( .ip1(n13253), .ip2(\cache_tag_B[3][6] ), .ip3(n9049), .ip4(n9048), .op(n9051) );
  nand2_1 U9239 ( .ip1(n13278), .ip2(\cache_tag_B[1][6] ), .op(n9050) );
  nand3_1 U9240 ( .ip1(n9052), .ip2(n9051), .ip3(n9050), .op(n9053) );
  xor2_1 U9241 ( .ip1(addr_req[13]), .ip2(n9053), .op(n9090) );
  nand2_1 U9242 ( .ip1(n9271), .ip2(\cache_tag_B[3][4] ), .op(n9063) );
  nor2_1 U9243 ( .ip1(n9178), .ip2(n9054), .op(n9060) );
  nand2_1 U9244 ( .ip1(n13268), .ip2(\cache_tag_B[4][4] ), .op(n9058) );
  nand2_1 U9245 ( .ip1(n13270), .ip2(\cache_tag_B[0][4] ), .op(n9057) );
  nand2_1 U9246 ( .ip1(n13269), .ip2(\cache_tag_B[6][4] ), .op(n9056) );
  nand2_1 U9247 ( .ip1(n13278), .ip2(\cache_tag_B[1][4] ), .op(n9055) );
  nand4_1 U9248 ( .ip1(n9058), .ip2(n9057), .ip3(n9056), .ip4(n9055), .op(
        n9059) );
  not_ab_or_c_or_d U9249 ( .ip1(n13264), .ip2(\cache_tag_B[2][4] ), .ip3(n9060), .ip4(n9059), .op(n9062) );
  nand2_1 U9250 ( .ip1(n13254), .ip2(\cache_tag_B[5][4] ), .op(n9061) );
  nand3_1 U9251 ( .ip1(n9063), .ip2(n9062), .ip3(n9061), .op(n9064) );
  xor2_1 U9252 ( .ip1(addr_req[11]), .ip2(n9064), .op(n9089) );
  nand2_1 U9253 ( .ip1(n13268), .ip2(\cache_tag_B[4][19] ), .op(n9074) );
  inv_1 U9254 ( .ip(n13277), .op(n9178) );
  nor2_1 U9255 ( .ip1(n9178), .ip2(n9065), .op(n9071) );
  nand2_1 U9256 ( .ip1(n13264), .ip2(\cache_tag_B[2][19] ), .op(n9069) );
  nand2_1 U9257 ( .ip1(n13253), .ip2(\cache_tag_B[3][19] ), .op(n9068) );
  nand2_1 U9258 ( .ip1(n13269), .ip2(\cache_tag_B[6][19] ), .op(n9067) );
  nand2_1 U9259 ( .ip1(n13254), .ip2(\cache_tag_B[5][19] ), .op(n9066) );
  nand4_1 U9260 ( .ip1(n9069), .ip2(n9068), .ip3(n9067), .ip4(n9066), .op(
        n9070) );
  not_ab_or_c_or_d U9261 ( .ip1(n13270), .ip2(\cache_tag_B[0][19] ), .ip3(
        n9071), .ip4(n9070), .op(n9073) );
  nand2_1 U9262 ( .ip1(n13278), .ip2(\cache_tag_B[1][19] ), .op(n9072) );
  nand3_1 U9263 ( .ip1(n9074), .ip2(n9073), .ip3(n9072), .op(n9075) );
  xor2_1 U9264 ( .ip1(addr_req[26]), .ip2(n9075), .op(n9088) );
  nand2_1 U9265 ( .ip1(n13268), .ip2(\cache_tag_B[4][0] ), .op(n9085) );
  nor2_1 U9266 ( .ip1(n9178), .ip2(n9076), .op(n9082) );
  nand2_1 U9267 ( .ip1(n13269), .ip2(\cache_tag_B[6][0] ), .op(n9080) );
  nand2_1 U9268 ( .ip1(n13278), .ip2(\cache_tag_B[1][0] ), .op(n9079) );
  nand2_1 U9269 ( .ip1(n13267), .ip2(\cache_tag_B[5][0] ), .op(n9078) );
  nand2_1 U9270 ( .ip1(n13270), .ip2(\cache_tag_B[0][0] ), .op(n9077) );
  nand4_1 U9271 ( .ip1(n9080), .ip2(n9079), .ip3(n9078), .ip4(n9077), .op(
        n9081) );
  not_ab_or_c_or_d U9272 ( .ip1(n13253), .ip2(\cache_tag_B[3][0] ), .ip3(n9082), .ip4(n9081), .op(n9084) );
  nand2_1 U9273 ( .ip1(n13264), .ip2(\cache_tag_B[2][0] ), .op(n9083) );
  nand3_1 U9274 ( .ip1(n9085), .ip2(n9084), .ip3(n9083), .op(n9086) );
  xor2_1 U9275 ( .ip1(addr_req[7]), .ip2(n9086), .op(n9087) );
  nor4_1 U9276 ( .ip1(n9090), .ip2(n9089), .ip3(n9088), .ip4(n9087), .op(n9317) );
  nand2_1 U9277 ( .ip1(\cache_tag_B[6][17] ), .ip2(n13251), .op(n9100) );
  nor2_1 U9278 ( .ip1(n9178), .ip2(n9091), .op(n9097) );
  nand2_1 U9279 ( .ip1(n13254), .ip2(\cache_tag_B[5][17] ), .op(n9095) );
  nand2_1 U9280 ( .ip1(n13278), .ip2(\cache_tag_B[1][17] ), .op(n9094) );
  nand2_1 U9281 ( .ip1(n13268), .ip2(\cache_tag_B[4][17] ), .op(n9093) );
  nand2_1 U9282 ( .ip1(n13264), .ip2(\cache_tag_B[2][17] ), .op(n9092) );
  nand4_1 U9283 ( .ip1(n9095), .ip2(n9094), .ip3(n9093), .ip4(n9092), .op(
        n9096) );
  not_ab_or_c_or_d U9284 ( .ip1(n9271), .ip2(\cache_tag_B[3][17] ), .ip3(n9097), .ip4(n9096), .op(n9099) );
  nand2_1 U9285 ( .ip1(n13270), .ip2(\cache_tag_B[0][17] ), .op(n9098) );
  nand3_1 U9286 ( .ip1(n9100), .ip2(n9099), .ip3(n9098), .op(n9101) );
  xor2_1 U9287 ( .ip1(addr_req[24]), .ip2(n9101), .op(n9139) );
  nand2_1 U9288 ( .ip1(\cache_tag_B[4][16] ), .ip2(n9102), .op(n9112) );
  nor2_1 U9289 ( .ip1(n9178), .ip2(n9103), .op(n9109) );
  nand2_1 U9290 ( .ip1(n13269), .ip2(\cache_tag_B[6][16] ), .op(n9107) );
  nand2_1 U9291 ( .ip1(n13253), .ip2(\cache_tag_B[3][16] ), .op(n9106) );
  nand2_1 U9292 ( .ip1(n13264), .ip2(\cache_tag_B[2][16] ), .op(n9105) );
  nand2_1 U9293 ( .ip1(n13267), .ip2(\cache_tag_B[5][16] ), .op(n9104) );
  nand4_1 U9294 ( .ip1(n9107), .ip2(n9106), .ip3(n9105), .ip4(n9104), .op(
        n9108) );
  not_ab_or_c_or_d U9295 ( .ip1(\cache_tag_B[0][16] ), .ip2(n13270), .ip3(
        n9109), .ip4(n9108), .op(n9111) );
  nand2_1 U9296 ( .ip1(n13278), .ip2(\cache_tag_B[1][16] ), .op(n9110) );
  nand3_1 U9297 ( .ip1(n9112), .ip2(n9111), .ip3(n9110), .op(n9113) );
  xor2_1 U9298 ( .ip1(addr_req[23]), .ip2(n9113), .op(n9138) );
  nand2_1 U9299 ( .ip1(n13269), .ip2(\cache_tag_B[6][9] ), .op(n9123) );
  nor2_1 U9300 ( .ip1(n9178), .ip2(n9114), .op(n9120) );
  nand2_1 U9301 ( .ip1(n13268), .ip2(\cache_tag_B[4][9] ), .op(n9118) );
  nand2_1 U9302 ( .ip1(n13278), .ip2(\cache_tag_B[1][9] ), .op(n9117) );
  nand2_1 U9303 ( .ip1(n13264), .ip2(\cache_tag_B[2][9] ), .op(n9116) );
  nand2_1 U9304 ( .ip1(n13253), .ip2(\cache_tag_B[3][9] ), .op(n9115) );
  nand4_1 U9305 ( .ip1(n9118), .ip2(n9117), .ip3(n9116), .ip4(n9115), .op(
        n9119) );
  not_ab_or_c_or_d U9306 ( .ip1(n13270), .ip2(\cache_tag_B[0][9] ), .ip3(n9120), .ip4(n9119), .op(n9122) );
  nand2_1 U9307 ( .ip1(n13267), .ip2(\cache_tag_B[5][9] ), .op(n9121) );
  nand3_1 U9308 ( .ip1(n9123), .ip2(n9122), .ip3(n9121), .op(n9124) );
  xor2_1 U9309 ( .ip1(addr_req[16]), .ip2(n9124), .op(n9137) );
  nand2_1 U9310 ( .ip1(\cache_tag_B[3][8] ), .ip2(n13253), .op(n9134) );
  nor2_1 U9311 ( .ip1(n9178), .ip2(n9125), .op(n9131) );
  nand2_1 U9312 ( .ip1(n13278), .ip2(\cache_tag_B[1][8] ), .op(n9129) );
  nand2_1 U9313 ( .ip1(n13269), .ip2(\cache_tag_B[6][8] ), .op(n9128) );
  nand2_1 U9314 ( .ip1(n13268), .ip2(\cache_tag_B[4][8] ), .op(n9127) );
  nand2_1 U9315 ( .ip1(n13270), .ip2(\cache_tag_B[0][8] ), .op(n9126) );
  nand4_1 U9316 ( .ip1(n9129), .ip2(n9128), .ip3(n9127), .ip4(n9126), .op(
        n9130) );
  not_ab_or_c_or_d U9317 ( .ip1(n13264), .ip2(\cache_tag_B[2][8] ), .ip3(n9131), .ip4(n9130), .op(n9133) );
  nand2_1 U9318 ( .ip1(n13254), .ip2(\cache_tag_B[5][8] ), .op(n9132) );
  nand3_1 U9319 ( .ip1(n9134), .ip2(n9133), .ip3(n9132), .op(n9135) );
  xor2_1 U9320 ( .ip1(addr_req[15]), .ip2(n9135), .op(n9136) );
  nor4_1 U9321 ( .ip1(n9139), .ip2(n9138), .ip3(n9137), .ip4(n9136), .op(n9316) );
  nand2_1 U9322 ( .ip1(\cache_tag_B[0][24] ), .ip2(n13270), .op(n9149) );
  nor2_1 U9323 ( .ip1(n9178), .ip2(n9140), .op(n9146) );
  nand2_1 U9324 ( .ip1(n13264), .ip2(\cache_tag_B[2][24] ), .op(n9144) );
  nand2_1 U9325 ( .ip1(n13278), .ip2(\cache_tag_B[1][24] ), .op(n9143) );
  nand2_1 U9326 ( .ip1(n13268), .ip2(\cache_tag_B[4][24] ), .op(n9142) );
  nand2_1 U9327 ( .ip1(n13267), .ip2(\cache_tag_B[5][24] ), .op(n9141) );
  nand4_1 U9328 ( .ip1(n9144), .ip2(n9143), .ip3(n9142), .ip4(n9141), .op(
        n9145) );
  not_ab_or_c_or_d U9329 ( .ip1(\cache_tag_B[6][24] ), .ip2(n13251), .ip3(
        n9146), .ip4(n9145), .op(n9148) );
  nand2_1 U9330 ( .ip1(n13253), .ip2(\cache_tag_B[3][24] ), .op(n9147) );
  nand3_1 U9331 ( .ip1(n9149), .ip2(n9148), .ip3(n9147), .op(n9150) );
  xor2_1 U9332 ( .ip1(addr_req[31]), .ip2(n9150), .op(n9314) );
  nand2_1 U9333 ( .ip1(\cache_tag_B[2][1] ), .ip2(n9349), .op(n9160) );
  nor2_1 U9334 ( .ip1(n9178), .ip2(n9151), .op(n9157) );
  nand2_1 U9335 ( .ip1(n13268), .ip2(\cache_tag_B[4][1] ), .op(n9155) );
  nand2_1 U9336 ( .ip1(n13253), .ip2(\cache_tag_B[3][1] ), .op(n9154) );
  nand2_1 U9337 ( .ip1(n13269), .ip2(\cache_tag_B[6][1] ), .op(n9153) );
  nand2_1 U9338 ( .ip1(n13267), .ip2(\cache_tag_B[5][1] ), .op(n9152) );
  nand4_1 U9339 ( .ip1(n9155), .ip2(n9154), .ip3(n9153), .ip4(n9152), .op(
        n9156) );
  not_ab_or_c_or_d U9340 ( .ip1(\cache_tag_B[1][1] ), .ip2(n13278), .ip3(n9157), .ip4(n9156), .op(n9159) );
  nand2_1 U9341 ( .ip1(n13270), .ip2(\cache_tag_B[0][1] ), .op(n9158) );
  nand3_1 U9342 ( .ip1(n9160), .ip2(n9159), .ip3(n9158), .op(n9161) );
  mux2_1 U9343 ( .ip1(n9162), .ip2(addr_req[8]), .s(n9161), .op(n9205) );
  inv_1 U9344 ( .ip(addr_req[21]), .op(n9176) );
  nand2_1 U9345 ( .ip1(\cache_tag_B[6][14] ), .ip2(n13251), .op(n9174) );
  nor2_1 U9346 ( .ip1(n9164), .ip2(n9163), .op(n9171) );
  nand2_1 U9347 ( .ip1(n13277), .ip2(\cache_tag_B[7][14] ), .op(n9169) );
  nand2_1 U9348 ( .ip1(n13268), .ip2(\cache_tag_B[4][14] ), .op(n9168) );
  nand2_1 U9349 ( .ip1(n9165), .ip2(\cache_tag_B[0][14] ), .op(n9167) );
  nand2_1 U9350 ( .ip1(n13278), .ip2(\cache_tag_B[1][14] ), .op(n9166) );
  nand4_1 U9351 ( .ip1(n9169), .ip2(n9168), .ip3(n9167), .ip4(n9166), .op(
        n9170) );
  not_ab_or_c_or_d U9352 ( .ip1(n13264), .ip2(\cache_tag_B[2][14] ), .ip3(
        n9171), .ip4(n9170), .op(n9173) );
  nand2_1 U9353 ( .ip1(n9271), .ip2(\cache_tag_B[3][14] ), .op(n9172) );
  nand3_1 U9354 ( .ip1(n9174), .ip2(n9173), .ip3(n9172), .op(n9175) );
  mux2_1 U9355 ( .ip1(n9176), .ip2(addr_req[21]), .s(n9175), .op(n9204) );
  nand2_1 U9356 ( .ip1(n13253), .ip2(\cache_tag_B[3][12] ), .op(n9187) );
  nor2_1 U9357 ( .ip1(n9178), .ip2(n9177), .op(n9184) );
  nand2_1 U9358 ( .ip1(n13264), .ip2(\cache_tag_B[2][12] ), .op(n9182) );
  nand2_1 U9359 ( .ip1(n13267), .ip2(\cache_tag_B[5][12] ), .op(n9181) );
  nand2_1 U9360 ( .ip1(n13278), .ip2(\cache_tag_B[1][12] ), .op(n9180) );
  nand2_1 U9361 ( .ip1(n13269), .ip2(\cache_tag_B[6][12] ), .op(n9179) );
  nand4_1 U9362 ( .ip1(n9182), .ip2(n9181), .ip3(n9180), .ip4(n9179), .op(
        n9183) );
  not_ab_or_c_or_d U9363 ( .ip1(n13268), .ip2(\cache_tag_B[4][12] ), .ip3(
        n9184), .ip4(n9183), .op(n9186) );
  nand2_1 U9364 ( .ip1(n13270), .ip2(\cache_tag_B[0][12] ), .op(n9185) );
  nand3_1 U9365 ( .ip1(n9187), .ip2(n9186), .ip3(n9185), .op(n9188) );
  mux2_1 U9366 ( .ip1(n9189), .ip2(addr_req[19]), .s(n9188), .op(n9203) );
  inv_1 U9367 ( .ip(addr_req[18]), .op(n9201) );
  nand2_1 U9368 ( .ip1(\cache_tag_B[3][11] ), .ip2(n13253), .op(n9199) );
  nor2_1 U9369 ( .ip1(n9178), .ip2(n9190), .op(n9196) );
  nand2_1 U9370 ( .ip1(n13267), .ip2(\cache_tag_B[5][11] ), .op(n9194) );
  nand2_1 U9371 ( .ip1(n13278), .ip2(\cache_tag_B[1][11] ), .op(n9193) );
  nand2_1 U9372 ( .ip1(n13269), .ip2(\cache_tag_B[6][11] ), .op(n9192) );
  nand2_1 U9373 ( .ip1(n13264), .ip2(\cache_tag_B[2][11] ), .op(n9191) );
  nand4_1 U9374 ( .ip1(n9194), .ip2(n9193), .ip3(n9192), .ip4(n9191), .op(
        n9195) );
  not_ab_or_c_or_d U9375 ( .ip1(n13268), .ip2(\cache_tag_B[4][11] ), .ip3(
        n9196), .ip4(n9195), .op(n9198) );
  nand2_1 U9376 ( .ip1(n13270), .ip2(\cache_tag_B[0][11] ), .op(n9197) );
  nand3_1 U9377 ( .ip1(n9199), .ip2(n9198), .ip3(n9197), .op(n9200) );
  mux2_1 U9378 ( .ip1(n9201), .ip2(addr_req[18]), .s(n9200), .op(n9202) );
  nand4_1 U9379 ( .ip1(n9205), .ip2(n9204), .ip3(n9203), .ip4(n9202), .op(
        n9313) );
  nand2_1 U9380 ( .ip1(n13267), .ip2(\cache_tag_B[5][15] ), .op(n9215) );
  nor2_1 U9381 ( .ip1(n9178), .ip2(n9206), .op(n9212) );
  nand2_1 U9382 ( .ip1(n9349), .ip2(\cache_tag_B[2][15] ), .op(n9210) );
  nand2_1 U9383 ( .ip1(n13270), .ip2(\cache_tag_B[0][15] ), .op(n9209) );
  nand2_1 U9384 ( .ip1(n13269), .ip2(\cache_tag_B[6][15] ), .op(n9208) );
  nand2_1 U9385 ( .ip1(n13253), .ip2(\cache_tag_B[3][15] ), .op(n9207) );
  nand4_1 U9386 ( .ip1(n9210), .ip2(n9209), .ip3(n9208), .ip4(n9207), .op(
        n9211) );
  not_ab_or_c_or_d U9387 ( .ip1(\cache_tag_B[4][15] ), .ip2(n13268), .ip3(
        n9212), .ip4(n9211), .op(n9214) );
  nand2_1 U9388 ( .ip1(n9225), .ip2(\cache_tag_B[1][15] ), .op(n9213) );
  nand3_1 U9389 ( .ip1(n9215), .ip2(n9214), .ip3(n9213), .op(n9216) );
  mux2_1 U9390 ( .ip1(n9217), .ip2(addr_req[22]), .s(n9216), .op(n9257) );
  inv_1 U9391 ( .ip(addr_req[9]), .op(n9230) );
  nand2_1 U9392 ( .ip1(n9349), .ip2(\cache_tag_B[2][2] ), .op(n9228) );
  nor2_1 U9393 ( .ip1(n13266), .ip2(n9218), .op(n9224) );
  nand2_1 U9394 ( .ip1(n13269), .ip2(\cache_tag_B[6][2] ), .op(n9222) );
  nand2_1 U9395 ( .ip1(n13268), .ip2(\cache_tag_B[4][2] ), .op(n9221) );
  nand2_1 U9396 ( .ip1(n13254), .ip2(\cache_tag_B[5][2] ), .op(n9220) );
  nand2_1 U9397 ( .ip1(n13277), .ip2(\cache_tag_B[7][2] ), .op(n9219) );
  nand4_1 U9398 ( .ip1(n9222), .ip2(n9221), .ip3(n9220), .ip4(n9219), .op(
        n9223) );
  not_ab_or_c_or_d U9399 ( .ip1(\cache_tag_B[1][2] ), .ip2(n9225), .ip3(n9224), 
        .ip4(n9223), .op(n9227) );
  nand2_1 U9400 ( .ip1(n13270), .ip2(\cache_tag_B[0][2] ), .op(n9226) );
  nand3_1 U9401 ( .ip1(n9228), .ip2(n9227), .ip3(n9226), .op(n9229) );
  mux2_1 U9402 ( .ip1(n9230), .ip2(addr_req[9]), .s(n9229), .op(n9256) );
  inv_1 U9403 ( .ip(addr_req[14]), .op(n9241) );
  nand2_1 U9404 ( .ip1(\cache_tag_B[4][7] ), .ip2(n13268), .op(n9239) );
  and2_1 U9405 ( .ip1(n13264), .ip2(\cache_tag_B[2][7] ), .op(n9236) );
  nand2_1 U9406 ( .ip1(n13277), .ip2(\cache_tag_B[7][7] ), .op(n9234) );
  nand2_1 U9407 ( .ip1(n13253), .ip2(\cache_tag_B[3][7] ), .op(n9233) );
  nand2_1 U9408 ( .ip1(n13267), .ip2(\cache_tag_B[5][7] ), .op(n9232) );
  nand2_1 U9409 ( .ip1(n13278), .ip2(\cache_tag_B[1][7] ), .op(n9231) );
  nand4_1 U9410 ( .ip1(n9234), .ip2(n9233), .ip3(n9232), .ip4(n9231), .op(
        n9235) );
  not_ab_or_c_or_d U9411 ( .ip1(\cache_tag_B[6][7] ), .ip2(n13251), .ip3(n9236), .ip4(n9235), .op(n9238) );
  nand2_1 U9412 ( .ip1(n13270), .ip2(\cache_tag_B[0][7] ), .op(n9237) );
  nand3_1 U9413 ( .ip1(n9239), .ip2(n9238), .ip3(n9237), .op(n9240) );
  mux2_1 U9414 ( .ip1(n9241), .ip2(addr_req[14]), .s(n9240), .op(n9255) );
  inv_1 U9415 ( .ip(addr_req[30]), .op(n9253) );
  nand2_1 U9416 ( .ip1(\cache_tag_B[2][23] ), .ip2(n9349), .op(n9251) );
  nor2_1 U9417 ( .ip1(n13266), .ip2(n9242), .op(n9248) );
  nand2_1 U9418 ( .ip1(n13268), .ip2(\cache_tag_B[4][23] ), .op(n9246) );
  nand2_1 U9419 ( .ip1(n13269), .ip2(\cache_tag_B[6][23] ), .op(n9245) );
  nand2_1 U9420 ( .ip1(n13254), .ip2(\cache_tag_B[5][23] ), .op(n9244) );
  nand2_1 U9421 ( .ip1(n13277), .ip2(\cache_tag_B[7][23] ), .op(n9243) );
  nand4_1 U9422 ( .ip1(n9246), .ip2(n9245), .ip3(n9244), .ip4(n9243), .op(
        n9247) );
  not_ab_or_c_or_d U9423 ( .ip1(n13278), .ip2(\cache_tag_B[1][23] ), .ip3(
        n9248), .ip4(n9247), .op(n9250) );
  nand2_1 U9424 ( .ip1(n13270), .ip2(\cache_tag_B[0][23] ), .op(n9249) );
  nand3_1 U9425 ( .ip1(n9251), .ip2(n9250), .ip3(n9249), .op(n9252) );
  mux2_1 U9426 ( .ip1(n9253), .ip2(addr_req[30]), .s(n9252), .op(n9254) );
  nand4_1 U9427 ( .ip1(n9257), .ip2(n9256), .ip3(n9255), .ip4(n9254), .op(
        n9312) );
  inv_1 U9428 ( .ip(addr_req[20]), .op(n9269) );
  nand2_1 U9429 ( .ip1(n13253), .ip2(\cache_tag_B[3][13] ), .op(n9267) );
  nor2_1 U9430 ( .ip1(n9178), .ip2(n9258), .op(n9264) );
  nand2_1 U9431 ( .ip1(n13270), .ip2(\cache_tag_B[0][13] ), .op(n9262) );
  nand2_1 U9432 ( .ip1(n13264), .ip2(\cache_tag_B[2][13] ), .op(n9261) );
  nand2_1 U9433 ( .ip1(n13268), .ip2(\cache_tag_B[4][13] ), .op(n9260) );
  nand2_1 U9434 ( .ip1(n13254), .ip2(\cache_tag_B[5][13] ), .op(n9259) );
  nand4_1 U9435 ( .ip1(n9262), .ip2(n9261), .ip3(n9260), .ip4(n9259), .op(
        n9263) );
  not_ab_or_c_or_d U9436 ( .ip1(\cache_tag_B[6][13] ), .ip2(n13251), .ip3(
        n9264), .ip4(n9263), .op(n9266) );
  nand2_1 U9437 ( .ip1(n13278), .ip2(\cache_tag_B[1][13] ), .op(n9265) );
  nand3_1 U9438 ( .ip1(n9267), .ip2(n9266), .ip3(n9265), .op(n9268) );
  mux2_1 U9439 ( .ip1(n9269), .ip2(addr_req[20]), .s(n9268), .op(n9310) );
  inv_1 U9440 ( .ip(addr_req[28]), .op(n9282) );
  nand2_1 U9441 ( .ip1(\cache_tag_B[6][21] ), .ip2(n13251), .op(n9280) );
  nor2_1 U9442 ( .ip1(n9178), .ip2(n9270), .op(n9277) );
  nand2_1 U9443 ( .ip1(n13278), .ip2(\cache_tag_B[1][21] ), .op(n9275) );
  nand2_1 U9444 ( .ip1(n13268), .ip2(\cache_tag_B[4][21] ), .op(n9274) );
  nand2_1 U9445 ( .ip1(n13254), .ip2(\cache_tag_B[5][21] ), .op(n9273) );
  nand2_1 U9446 ( .ip1(n9271), .ip2(\cache_tag_B[3][21] ), .op(n9272) );
  nand4_1 U9447 ( .ip1(n9275), .ip2(n9274), .ip3(n9273), .ip4(n9272), .op(
        n9276) );
  not_ab_or_c_or_d U9448 ( .ip1(\cache_tag_B[2][21] ), .ip2(n9349), .ip3(n9277), .ip4(n9276), .op(n9279) );
  nand2_1 U9449 ( .ip1(n13270), .ip2(\cache_tag_B[0][21] ), .op(n9278) );
  nand3_1 U9450 ( .ip1(n9280), .ip2(n9279), .ip3(n9278), .op(n9281) );
  mux2_1 U9451 ( .ip1(n9282), .ip2(addr_req[28]), .s(n9281), .op(n9309) );
  inv_1 U9452 ( .ip(addr_req[17]), .op(n9294) );
  nand2_1 U9453 ( .ip1(n9349), .ip2(\cache_tag_B[2][10] ), .op(n9292) );
  nor2_1 U9454 ( .ip1(n9178), .ip2(n9283), .op(n9289) );
  nand2_1 U9455 ( .ip1(n13269), .ip2(\cache_tag_B[6][10] ), .op(n9287) );
  nand2_1 U9456 ( .ip1(n13253), .ip2(\cache_tag_B[3][10] ), .op(n9286) );
  nand2_1 U9457 ( .ip1(n13278), .ip2(\cache_tag_B[1][10] ), .op(n9285) );
  nand2_1 U9458 ( .ip1(n13270), .ip2(\cache_tag_B[0][10] ), .op(n9284) );
  nand4_1 U9459 ( .ip1(n9287), .ip2(n9286), .ip3(n9285), .ip4(n9284), .op(
        n9288) );
  not_ab_or_c_or_d U9460 ( .ip1(\cache_tag_B[4][10] ), .ip2(n13268), .ip3(
        n9289), .ip4(n9288), .op(n9291) );
  nand2_1 U9461 ( .ip1(n13254), .ip2(\cache_tag_B[5][10] ), .op(n9290) );
  nand3_1 U9462 ( .ip1(n9292), .ip2(n9291), .ip3(n9290), .op(n9293) );
  mux2_1 U9463 ( .ip1(n9294), .ip2(addr_req[17]), .s(n9293), .op(n9308) );
  nand2_1 U9464 ( .ip1(\cache_tag_B[0][22] ), .ip2(n13270), .op(n9304) );
  nor2_1 U9465 ( .ip1(n9178), .ip2(n9295), .op(n9301) );
  nand2_1 U9466 ( .ip1(n13264), .ip2(\cache_tag_B[2][22] ), .op(n9299) );
  nand2_1 U9467 ( .ip1(n13251), .ip2(\cache_tag_B[6][22] ), .op(n9298) );
  nand2_1 U9468 ( .ip1(n13268), .ip2(\cache_tag_B[4][22] ), .op(n9297) );
  nand2_1 U9469 ( .ip1(n13254), .ip2(\cache_tag_B[5][22] ), .op(n9296) );
  nand4_1 U9470 ( .ip1(n9299), .ip2(n9298), .ip3(n9297), .ip4(n9296), .op(
        n9300) );
  not_ab_or_c_or_d U9471 ( .ip1(n13278), .ip2(\cache_tag_B[1][22] ), .ip3(
        n9301), .ip4(n9300), .op(n9303) );
  nand2_1 U9472 ( .ip1(n13253), .ip2(\cache_tag_B[3][22] ), .op(n9302) );
  nand3_1 U9473 ( .ip1(n9304), .ip2(n9303), .ip3(n9302), .op(n9305) );
  mux2_1 U9474 ( .ip1(n9306), .ip2(addr_req[29]), .s(n9305), .op(n9307) );
  nand4_1 U9475 ( .ip1(n9310), .ip2(n9309), .ip3(n9308), .ip4(n9307), .op(
        n9311) );
  nor4_1 U9476 ( .ip1(n9314), .ip2(n9313), .ip3(n9312), .ip4(n9311), .op(n9315) );
  nand4_1 U9477 ( .ip1(n9318), .ip2(n9317), .ip3(n9316), .ip4(n9315), .op(
        n13284) );
  inv_1 U9478 ( .ip(n13284), .op(n9319) );
  nor3_1 U9479 ( .ip1(n13290), .ip2(n13283), .ip3(n9319), .op(n9359) );
  nor2_1 U9480 ( .ip1(hit), .ip2(n9320), .op(n9321) );
  nor2_1 U9481 ( .ip1(n9359), .ip2(n9321), .op(n5188) );
  nand3_1 U9482 ( .ip1(n9324), .ip2(n9323), .ip3(n9322), .op(n9326) );
  nand2_1 U9483 ( .ip1(n9326), .ip2(n9325), .op(next_state[0]) );
  inv_1 U9484 ( .ip(next_state[0]), .op(N4447) );
  nand2_1 U9485 ( .ip1(n13251), .ip2(cache_dirty_A[6]), .op(n9335) );
  and2_1 U9486 ( .ip1(n13267), .ip2(cache_dirty_A[5]), .op(n9332) );
  nand2_1 U9487 ( .ip1(n13270), .ip2(cache_dirty_A[0]), .op(n9330) );
  nand2_1 U9488 ( .ip1(n13253), .ip2(cache_dirty_A[3]), .op(n9329) );
  nand2_1 U9489 ( .ip1(n13278), .ip2(cache_dirty_A[1]), .op(n9328) );
  nand2_1 U9490 ( .ip1(n13268), .ip2(cache_dirty_A[4]), .op(n9327) );
  nand4_1 U9491 ( .ip1(n9330), .ip2(n9329), .ip3(n9328), .ip4(n9327), .op(
        n9331) );
  not_ab_or_c_or_d U9492 ( .ip1(cache_dirty_A[7]), .ip2(n13277), .ip3(n9332), 
        .ip4(n9331), .op(n9334) );
  nand2_1 U9493 ( .ip1(n13264), .ip2(cache_dirty_A[2]), .op(n9333) );
  nand3_1 U9494 ( .ip1(n9335), .ip2(n9334), .ip3(n9333), .op(n9357) );
  nand2_1 U9495 ( .ip1(n13254), .ip2(cache_dirty_B[5]), .op(n9344) );
  and2_1 U9496 ( .ip1(n13251), .ip2(cache_dirty_B[6]), .op(n9341) );
  nand2_1 U9497 ( .ip1(n13253), .ip2(cache_dirty_B[3]), .op(n9339) );
  nand2_1 U9498 ( .ip1(n13277), .ip2(cache_dirty_B[7]), .op(n9338) );
  nand2_1 U9499 ( .ip1(n13268), .ip2(cache_dirty_B[4]), .op(n9337) );
  nand2_1 U9500 ( .ip1(n13264), .ip2(cache_dirty_B[2]), .op(n9336) );
  nand4_1 U9501 ( .ip1(n9339), .ip2(n9338), .ip3(n9337), .ip4(n9336), .op(
        n9340) );
  not_ab_or_c_or_d U9502 ( .ip1(cache_dirty_B[0]), .ip2(n13270), .ip3(n9341), 
        .ip4(n9340), .op(n9343) );
  nand2_1 U9503 ( .ip1(n13278), .ip2(cache_dirty_B[1]), .op(n9342) );
  nand3_1 U9504 ( .ip1(n9344), .ip2(n9343), .ip3(n9342), .op(n9356) );
  nand2_1 U9505 ( .ip1(n13254), .ip2(cache_line_count[5]), .op(n9348) );
  nand2_1 U9506 ( .ip1(n13270), .ip2(cache_line_count[0]), .op(n9347) );
  nand2_1 U9507 ( .ip1(n13268), .ip2(cache_line_count[4]), .op(n9346) );
  nand2_1 U9508 ( .ip1(n13277), .ip2(cache_line_count[7]), .op(n9345) );
  nand4_1 U9509 ( .ip1(n9348), .ip2(n9347), .ip3(n9346), .ip4(n9345), .op(
        n9355) );
  nand2_1 U9510 ( .ip1(n9349), .ip2(cache_line_count[2]), .op(n9353) );
  nand2_1 U9511 ( .ip1(n13278), .ip2(cache_line_count[1]), .op(n9352) );
  nand2_1 U9512 ( .ip1(n13251), .ip2(cache_line_count[6]), .op(n9351) );
  nand2_1 U9513 ( .ip1(n13253), .ip2(cache_line_count[3]), .op(n9350) );
  nand4_1 U9514 ( .ip1(n9353), .ip2(n9352), .ip3(n9351), .ip4(n9350), .op(
        n9354) );
  nor2_1 U9515 ( .ip1(n9355), .ip2(n9354), .op(n13282) );
  inv_1 U9516 ( .ip(n13282), .op(n9361) );
  mux2_1 U9517 ( .ip1(n9357), .ip2(n9356), .s(n9361), .op(n9358) );
  mux2_1 U9518 ( .ip1(dirty), .ip2(n9358), .s(n9359), .op(n7941) );
  inv_1 U9519 ( .ip(n9359), .op(n13205) );
  nor2_1 U9520 ( .ip1(rst), .ip2(n13205), .op(n9360) );
  mux2_1 U9521 ( .ip1(SelectWay), .ip2(n9361), .s(n9360), .op(n7940) );
  or2_1 U9522 ( .ip1(n9363), .ip2(n9362), .op(n9407) );
  buf_1 U9523 ( .ip(n9407), .op(n9425) );
  nand2_1 U9524 ( .ip1(rd_temp), .ip2(n9425), .op(n9365) );
  nand2_1 U9525 ( .ip1(rd), .ip2(next_state[1]), .op(n9364) );
  nand2_1 U9526 ( .ip1(n9365), .ip2(n9364), .op(n7939) );
  mux2_1 U9527 ( .ip1(addr_req[0]), .ip2(N4300), .s(n9407), .op(n7938) );
  and2_1 U9528 ( .ip1(n9425), .ip2(N4301), .op(n7937) );
  mux2_1 U9529 ( .ip1(addr_req[1]), .ip2(N4297), .s(n9407), .op(n7936) );
  and2_1 U9530 ( .ip1(n9425), .ip2(N4298), .op(n7935) );
  mux2_1 U9531 ( .ip1(addr_req[2]), .ip2(N4294), .s(n9407), .op(n7934) );
  and2_1 U9532 ( .ip1(n9425), .ip2(N4295), .op(n7933) );
  mux2_1 U9533 ( .ip1(addr_req[3]), .ip2(N4291), .s(n9407), .op(n7932) );
  and2_1 U9534 ( .ip1(n9425), .ip2(N4292), .op(n7931) );
  mux2_1 U9535 ( .ip1(addr_req[4]), .ip2(N4288), .s(n9407), .op(n7930) );
  and2_1 U9536 ( .ip1(n9425), .ip2(N4289), .op(n7929) );
  mux2_1 U9537 ( .ip1(addr_req[5]), .ip2(N4285), .s(n9407), .op(n7928) );
  and2_1 U9538 ( .ip1(n9425), .ip2(N4286), .op(n7927) );
  mux2_1 U9539 ( .ip1(addr_req[6]), .ip2(N4282), .s(n9407), .op(n7926) );
  and2_1 U9540 ( .ip1(n9425), .ip2(N4283), .op(n7925) );
  nor2_1 U9541 ( .ip1(n12618), .ip2(n9860), .op(n9708) );
  nand2_1 U9542 ( .ip1(n9703), .ip2(n9708), .op(n9366) );
  mux2_1 U9543 ( .ip1(n9702), .ip2(cache_line_count[0]), .s(n9366), .op(n7924)
         );
  nor2_1 U9544 ( .ip1(n12618), .ip2(n9862), .op(n9717) );
  nand2_1 U9545 ( .ip1(n9703), .ip2(n9717), .op(n9367) );
  mux2_1 U9546 ( .ip1(n9702), .ip2(cache_line_count[1]), .s(n9367), .op(n7923)
         );
  nor2_1 U9547 ( .ip1(n12618), .ip2(n9864), .op(n9726) );
  nand2_1 U9548 ( .ip1(n9703), .ip2(n9726), .op(n9368) );
  mux2_1 U9549 ( .ip1(n9702), .ip2(cache_line_count[2]), .s(n9368), .op(n7922)
         );
  nor2_1 U9550 ( .ip1(rst), .ip2(n9866), .op(n9735) );
  nand2_1 U9551 ( .ip1(n9703), .ip2(n9735), .op(n9369) );
  mux2_1 U9552 ( .ip1(n9702), .ip2(cache_line_count[3]), .s(n9369), .op(n7921)
         );
  nor2_1 U9553 ( .ip1(n12618), .ip2(n9868), .op(n9744) );
  nand2_1 U9554 ( .ip1(n9703), .ip2(n9744), .op(n9370) );
  mux2_1 U9555 ( .ip1(n9702), .ip2(cache_line_count[4]), .s(n9370), .op(n7920)
         );
  nor2_1 U9556 ( .ip1(n12618), .ip2(n9870), .op(n9753) );
  nand2_1 U9557 ( .ip1(n9703), .ip2(n9753), .op(n9371) );
  mux2_1 U9558 ( .ip1(n9702), .ip2(cache_line_count[5]), .s(n9371), .op(n7919)
         );
  nor2_1 U9559 ( .ip1(n12618), .ip2(n9762), .op(n9765) );
  nand2_1 U9560 ( .ip1(n9703), .ip2(n9765), .op(n9372) );
  mux2_1 U9561 ( .ip1(n9702), .ip2(cache_line_count[6]), .s(n9372), .op(n7918)
         );
  nor2_1 U9562 ( .ip1(rst), .ip2(n9769), .op(n9811) );
  nand2_1 U9563 ( .ip1(n9703), .ip2(n9811), .op(n9373) );
  mux2_1 U9564 ( .ip1(n9702), .ip2(cache_line_count[7]), .s(n9373), .op(n7917)
         );
  nand2_1 U9565 ( .ip1(n9703), .ip2(SelectWay), .op(n9847) );
  nor2_1 U9566 ( .ip1(n9860), .ip2(n9847), .op(n9374) );
  or2_1 U9567 ( .ip1(cache_valid_B[0]), .ip2(n9374), .op(n7916) );
  nor2_1 U9568 ( .ip1(n9862), .ip2(n9847), .op(n9375) );
  or2_1 U9569 ( .ip1(cache_valid_B[1]), .ip2(n9375), .op(n7915) );
  nor2_1 U9570 ( .ip1(n9864), .ip2(n9847), .op(n9376) );
  or2_1 U9571 ( .ip1(cache_valid_B[2]), .ip2(n9376), .op(n7914) );
  inv_1 U9572 ( .ip(cache_valid_B[3]), .op(n13265) );
  or2_1 U9573 ( .ip1(n9866), .ip2(n9847), .op(n9377) );
  nand2_1 U9574 ( .ip1(n13265), .ip2(n9377), .op(n7913) );
  nor2_1 U9575 ( .ip1(n9868), .ip2(n9847), .op(n9378) );
  or2_1 U9576 ( .ip1(cache_valid_B[4]), .ip2(n9378), .op(n7912) );
  nor2_1 U9577 ( .ip1(n9870), .ip2(n9847), .op(n9379) );
  or2_1 U9578 ( .ip1(cache_valid_B[5]), .ip2(n9379), .op(n7911) );
  nor2_1 U9579 ( .ip1(n9762), .ip2(n9847), .op(n9380) );
  or2_1 U9580 ( .ip1(cache_valid_B[6]), .ip2(n9380), .op(n7910) );
  nor2_1 U9581 ( .ip1(n9769), .ip2(n9847), .op(n9381) );
  or2_1 U9582 ( .ip1(cache_valid_B[7]), .ip2(n9381), .op(n7909) );
  nand2_1 U9583 ( .ip1(n9702), .ip2(n9619), .op(n9389) );
  nor2_1 U9584 ( .ip1(n9860), .ip2(n9389), .op(n9382) );
  or2_1 U9585 ( .ip1(cache_valid_A[0]), .ip2(n9382), .op(n7908) );
  nor2_1 U9586 ( .ip1(n9862), .ip2(n9389), .op(n9383) );
  or2_1 U9587 ( .ip1(cache_valid_A[1]), .ip2(n9383), .op(n7907) );
  nor2_1 U9588 ( .ip1(n9864), .ip2(n9389), .op(n9384) );
  or2_1 U9589 ( .ip1(cache_valid_A[2]), .ip2(n9384), .op(n7906) );
  nor2_1 U9590 ( .ip1(n9866), .ip2(n9389), .op(n9385) );
  or2_1 U9591 ( .ip1(cache_valid_A[3]), .ip2(n9385), .op(n7905) );
  nor2_1 U9592 ( .ip1(n9868), .ip2(n9389), .op(n9386) );
  or2_1 U9593 ( .ip1(cache_valid_A[4]), .ip2(n9386), .op(n7904) );
  nor2_1 U9594 ( .ip1(n9870), .ip2(n9389), .op(n9387) );
  or2_1 U9595 ( .ip1(cache_valid_A[5]), .ip2(n9387), .op(n7903) );
  nor2_1 U9596 ( .ip1(n9762), .ip2(n9389), .op(n9388) );
  or2_1 U9597 ( .ip1(cache_valid_A[6]), .ip2(n9388), .op(n7902) );
  inv_1 U9598 ( .ip(cache_valid_A[7]), .op(n13252) );
  inv_1 U9599 ( .ip(n9389), .op(n9858) );
  nand2_1 U9600 ( .ip1(n10575), .ip2(n9858), .op(n9390) );
  nand2_1 U9601 ( .ip1(n13252), .ip2(n9390), .op(n7901) );
  mux2_1 U9602 ( .ip1(addr_req[7]), .ip2(N4279), .s(n9407), .op(n7900) );
  buf_1 U9603 ( .ip(n9407), .op(n9408) );
  and2_1 U9604 ( .ip1(n9408), .ip2(N4280), .op(n7899) );
  nand3_1 U9605 ( .ip1(n9703), .ip2(n9708), .ip3(n9702), .op(n9409) );
  buf_1 U9606 ( .ip(n9409), .op(n9391) );
  mux2_1 U9607 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[0][0] ), .s(n9391), 
        .op(n7898) );
  nand3_1 U9608 ( .ip1(n9703), .ip2(n9717), .ip3(n9702), .op(n9410) );
  buf_1 U9609 ( .ip(n9410), .op(n9392) );
  mux2_1 U9610 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[1][0] ), .s(n9392), 
        .op(n7897) );
  nand3_1 U9611 ( .ip1(n9703), .ip2(n9726), .ip3(n9702), .op(n9411) );
  buf_1 U9612 ( .ip(n9411), .op(n9393) );
  mux2_1 U9613 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[2][0] ), .s(n9393), 
        .op(n7896) );
  nand3_1 U9614 ( .ip1(n9619), .ip2(n9735), .ip3(n9702), .op(n9412) );
  buf_1 U9615 ( .ip(n9412), .op(n9394) );
  mux2_1 U9616 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[3][0] ), .s(n9394), 
        .op(n7895) );
  nand3_1 U9617 ( .ip1(n9703), .ip2(n9744), .ip3(n9702), .op(n9413) );
  buf_1 U9618 ( .ip(n9413), .op(n9395) );
  mux2_1 U9619 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[4][0] ), .s(n9395), 
        .op(n7894) );
  nand3_1 U9620 ( .ip1(n9703), .ip2(n9753), .ip3(n9702), .op(n9414) );
  buf_1 U9621 ( .ip(n9414), .op(n9396) );
  mux2_1 U9622 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[5][0] ), .s(n9396), 
        .op(n7893) );
  nand3_1 U9623 ( .ip1(n9703), .ip2(n9765), .ip3(n9702), .op(n9415) );
  buf_1 U9624 ( .ip(n9415), .op(n9397) );
  mux2_1 U9625 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[6][0] ), .s(n9397), 
        .op(n7892) );
  nand3_1 U9626 ( .ip1(n9703), .ip2(n9811), .ip3(n9702), .op(n9416) );
  buf_1 U9627 ( .ip(n9416), .op(n9398) );
  mux2_1 U9628 ( .ip1(addr_resp[7]), .ip2(\cache_tag_A[7][0] ), .s(n9398), 
        .op(n7891) );
  nand3_1 U9629 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9708), .op(n9417) );
  buf_1 U9630 ( .ip(n9417), .op(n9399) );
  mux2_1 U9631 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[0][0] ), .s(n9399), 
        .op(n7890) );
  nand3_1 U9632 ( .ip1(n9703), .ip2(SelectWay), .ip3(n9717), .op(n9418) );
  buf_1 U9633 ( .ip(n9418), .op(n9400) );
  mux2_1 U9634 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[1][0] ), .s(n9400), 
        .op(n7889) );
  nand3_1 U9635 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9726), .op(n9419) );
  buf_1 U9636 ( .ip(n9419), .op(n9401) );
  mux2_1 U9637 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[2][0] ), .s(n9401), 
        .op(n7888) );
  nand3_1 U9638 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9735), .op(n9420) );
  buf_1 U9639 ( .ip(n9420), .op(n9402) );
  mux2_1 U9640 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[3][0] ), .s(n9402), 
        .op(n7887) );
  nand3_1 U9641 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9744), .op(n9421) );
  buf_1 U9642 ( .ip(n9421), .op(n9403) );
  mux2_1 U9643 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[4][0] ), .s(n9403), 
        .op(n7886) );
  nand3_1 U9644 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9753), .op(n9422) );
  buf_1 U9645 ( .ip(n9422), .op(n9404) );
  mux2_1 U9646 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[5][0] ), .s(n9404), 
        .op(n7885) );
  nand3_1 U9647 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9765), .op(n9423) );
  buf_1 U9648 ( .ip(n9423), .op(n9405) );
  mux2_1 U9649 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[6][0] ), .s(n9405), 
        .op(n7884) );
  nand3_1 U9650 ( .ip1(n9619), .ip2(SelectWay), .ip3(n9811), .op(n9424) );
  buf_1 U9651 ( .ip(n9424), .op(n9406) );
  mux2_1 U9652 ( .ip1(addr_resp[7]), .ip2(\cache_tag_B[7][0] ), .s(n9406), 
        .op(n7883) );
  mux2_1 U9653 ( .ip1(addr_req[8]), .ip2(N4276), .s(n9408), .op(n7882) );
  and2_1 U9654 ( .ip1(n9425), .ip2(N4277), .op(n7881) );
  mux2_1 U9655 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[0][1] ), .s(n9391), 
        .op(n7880) );
  mux2_1 U9656 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[1][1] ), .s(n9392), 
        .op(n7879) );
  mux2_1 U9657 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[2][1] ), .s(n9393), 
        .op(n7878) );
  mux2_1 U9658 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[3][1] ), .s(n9394), 
        .op(n7877) );
  mux2_1 U9659 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[4][1] ), .s(n9395), 
        .op(n7876) );
  mux2_1 U9660 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[5][1] ), .s(n9396), 
        .op(n7875) );
  mux2_1 U9661 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[6][1] ), .s(n9397), 
        .op(n7874) );
  mux2_1 U9662 ( .ip1(addr_resp[8]), .ip2(\cache_tag_A[7][1] ), .s(n9398), 
        .op(n7873) );
  mux2_1 U9663 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[0][1] ), .s(n9399), 
        .op(n7872) );
  mux2_1 U9664 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[1][1] ), .s(n9400), 
        .op(n7871) );
  mux2_1 U9665 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[2][1] ), .s(n9401), 
        .op(n7870) );
  mux2_1 U9666 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[3][1] ), .s(n9402), 
        .op(n7869) );
  mux2_1 U9667 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[4][1] ), .s(n9403), 
        .op(n7868) );
  mux2_1 U9668 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[5][1] ), .s(n9404), 
        .op(n7867) );
  mux2_1 U9669 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[6][1] ), .s(n9405), 
        .op(n7866) );
  mux2_1 U9670 ( .ip1(addr_resp[8]), .ip2(\cache_tag_B[7][1] ), .s(n9406), 
        .op(n7865) );
  mux2_1 U9671 ( .ip1(addr_req[9]), .ip2(N4273), .s(n9408), .op(n7864) );
  and2_1 U9672 ( .ip1(n9425), .ip2(N4274), .op(n7863) );
  mux2_1 U9673 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[0][2] ), .s(n9391), 
        .op(n7862) );
  mux2_1 U9674 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[1][2] ), .s(n9392), 
        .op(n7861) );
  mux2_1 U9675 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[2][2] ), .s(n9393), 
        .op(n7860) );
  mux2_1 U9676 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[3][2] ), .s(n9394), 
        .op(n7859) );
  mux2_1 U9677 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[4][2] ), .s(n9395), 
        .op(n7858) );
  mux2_1 U9678 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[5][2] ), .s(n9396), 
        .op(n7857) );
  mux2_1 U9679 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[6][2] ), .s(n9397), 
        .op(n7856) );
  mux2_1 U9680 ( .ip1(addr_resp[9]), .ip2(\cache_tag_A[7][2] ), .s(n9398), 
        .op(n7855) );
  mux2_1 U9681 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[0][2] ), .s(n9399), 
        .op(n7854) );
  mux2_1 U9682 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[1][2] ), .s(n9400), 
        .op(n7853) );
  mux2_1 U9683 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[2][2] ), .s(n9401), 
        .op(n7852) );
  mux2_1 U9684 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[3][2] ), .s(n9402), 
        .op(n7851) );
  mux2_1 U9685 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[4][2] ), .s(n9403), 
        .op(n7850) );
  mux2_1 U9686 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[5][2] ), .s(n9404), 
        .op(n7849) );
  mux2_1 U9687 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[6][2] ), .s(n9405), 
        .op(n7848) );
  mux2_1 U9688 ( .ip1(addr_resp[9]), .ip2(\cache_tag_B[7][2] ), .s(n9406), 
        .op(n7847) );
  mux2_1 U9689 ( .ip1(addr_req[10]), .ip2(N4270), .s(n9408), .op(n7846) );
  and2_1 U9690 ( .ip1(n9425), .ip2(N4271), .op(n7845) );
  mux2_1 U9691 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[0][3] ), .s(n9391), 
        .op(n7844) );
  mux2_1 U9692 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[1][3] ), .s(n9392), 
        .op(n7843) );
  mux2_1 U9693 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[2][3] ), .s(n9393), 
        .op(n7842) );
  mux2_1 U9694 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[3][3] ), .s(n9394), 
        .op(n7841) );
  mux2_1 U9695 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[4][3] ), .s(n9395), 
        .op(n7840) );
  mux2_1 U9696 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[5][3] ), .s(n9396), 
        .op(n7839) );
  mux2_1 U9697 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[6][3] ), .s(n9397), 
        .op(n7838) );
  mux2_1 U9698 ( .ip1(addr_resp[10]), .ip2(\cache_tag_A[7][3] ), .s(n9398), 
        .op(n7837) );
  mux2_1 U9699 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[0][3] ), .s(n9399), 
        .op(n7836) );
  mux2_1 U9700 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[1][3] ), .s(n9400), 
        .op(n7835) );
  mux2_1 U9701 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[2][3] ), .s(n9401), 
        .op(n7834) );
  mux2_1 U9702 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[3][3] ), .s(n9402), 
        .op(n7833) );
  mux2_1 U9703 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[4][3] ), .s(n9403), 
        .op(n7832) );
  mux2_1 U9704 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[5][3] ), .s(n9404), 
        .op(n7831) );
  mux2_1 U9705 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[6][3] ), .s(n9405), 
        .op(n7830) );
  mux2_1 U9706 ( .ip1(addr_resp[10]), .ip2(\cache_tag_B[7][3] ), .s(n9406), 
        .op(n7829) );
  mux2_1 U9707 ( .ip1(addr_req[11]), .ip2(N4267), .s(n9407), .op(n7828) );
  and2_1 U9708 ( .ip1(n9425), .ip2(N4268), .op(n7827) );
  mux2_1 U9709 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[0][4] ), .s(n9391), 
        .op(n7826) );
  mux2_1 U9710 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[1][4] ), .s(n9392), 
        .op(n7825) );
  mux2_1 U9711 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[2][4] ), .s(n9393), 
        .op(n7824) );
  mux2_1 U9712 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[3][4] ), .s(n9394), 
        .op(n7823) );
  mux2_1 U9713 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[4][4] ), .s(n9395), 
        .op(n7822) );
  mux2_1 U9714 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[5][4] ), .s(n9396), 
        .op(n7821) );
  mux2_1 U9715 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[6][4] ), .s(n9397), 
        .op(n7820) );
  mux2_1 U9716 ( .ip1(addr_resp[11]), .ip2(\cache_tag_A[7][4] ), .s(n9398), 
        .op(n7819) );
  mux2_1 U9717 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[0][4] ), .s(n9399), 
        .op(n7818) );
  mux2_1 U9718 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[1][4] ), .s(n9400), 
        .op(n7817) );
  mux2_1 U9719 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[2][4] ), .s(n9401), 
        .op(n7816) );
  mux2_1 U9720 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[3][4] ), .s(n9402), 
        .op(n7815) );
  mux2_1 U9721 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[4][4] ), .s(n9403), 
        .op(n7814) );
  mux2_1 U9722 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[5][4] ), .s(n9404), 
        .op(n7813) );
  mux2_1 U9723 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[6][4] ), .s(n9405), 
        .op(n7812) );
  mux2_1 U9724 ( .ip1(addr_resp[11]), .ip2(\cache_tag_B[7][4] ), .s(n9406), 
        .op(n7811) );
  mux2_1 U9725 ( .ip1(addr_req[12]), .ip2(N4264), .s(n9408), .op(n7810) );
  and2_1 U9726 ( .ip1(n9425), .ip2(N4265), .op(n7809) );
  mux2_1 U9727 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[0][5] ), .s(n9391), 
        .op(n7808) );
  mux2_1 U9728 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[1][5] ), .s(n9392), 
        .op(n7807) );
  mux2_1 U9729 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[2][5] ), .s(n9393), 
        .op(n7806) );
  mux2_1 U9730 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[3][5] ), .s(n9394), 
        .op(n7805) );
  mux2_1 U9731 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[4][5] ), .s(n9395), 
        .op(n7804) );
  mux2_1 U9732 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[5][5] ), .s(n9396), 
        .op(n7803) );
  mux2_1 U9733 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[6][5] ), .s(n9397), 
        .op(n7802) );
  mux2_1 U9734 ( .ip1(addr_resp[12]), .ip2(\cache_tag_A[7][5] ), .s(n9398), 
        .op(n7801) );
  mux2_1 U9735 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[0][5] ), .s(n9399), 
        .op(n7800) );
  mux2_1 U9736 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[1][5] ), .s(n9400), 
        .op(n7799) );
  mux2_1 U9737 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[2][5] ), .s(n9401), 
        .op(n7798) );
  mux2_1 U9738 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[3][5] ), .s(n9402), 
        .op(n7797) );
  mux2_1 U9739 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[4][5] ), .s(n9403), 
        .op(n7796) );
  mux2_1 U9740 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[5][5] ), .s(n9404), 
        .op(n7795) );
  mux2_1 U9741 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[6][5] ), .s(n9405), 
        .op(n7794) );
  mux2_1 U9742 ( .ip1(addr_resp[12]), .ip2(\cache_tag_B[7][5] ), .s(n9406), 
        .op(n7793) );
  mux2_1 U9743 ( .ip1(addr_req[13]), .ip2(N4261), .s(n9408), .op(n7792) );
  and2_1 U9744 ( .ip1(n9425), .ip2(N4262), .op(n7791) );
  mux2_1 U9745 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[0][6] ), .s(n9391), 
        .op(n7790) );
  mux2_1 U9746 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[1][6] ), .s(n9392), 
        .op(n7789) );
  mux2_1 U9747 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[2][6] ), .s(n9393), 
        .op(n7788) );
  mux2_1 U9748 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[3][6] ), .s(n9394), 
        .op(n7787) );
  mux2_1 U9749 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[4][6] ), .s(n9395), 
        .op(n7786) );
  mux2_1 U9750 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[5][6] ), .s(n9396), 
        .op(n7785) );
  mux2_1 U9751 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[6][6] ), .s(n9397), 
        .op(n7784) );
  mux2_1 U9752 ( .ip1(addr_resp[13]), .ip2(\cache_tag_A[7][6] ), .s(n9398), 
        .op(n7783) );
  mux2_1 U9753 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[0][6] ), .s(n9399), 
        .op(n7782) );
  mux2_1 U9754 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[1][6] ), .s(n9400), 
        .op(n7781) );
  mux2_1 U9755 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[2][6] ), .s(n9401), 
        .op(n7780) );
  mux2_1 U9756 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[3][6] ), .s(n9402), 
        .op(n7779) );
  mux2_1 U9757 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[4][6] ), .s(n9403), 
        .op(n7778) );
  mux2_1 U9758 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[5][6] ), .s(n9404), 
        .op(n7777) );
  mux2_1 U9759 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[6][6] ), .s(n9405), 
        .op(n7776) );
  mux2_1 U9760 ( .ip1(addr_resp[13]), .ip2(\cache_tag_B[7][6] ), .s(n9406), 
        .op(n7775) );
  mux2_1 U9761 ( .ip1(addr_req[14]), .ip2(N4258), .s(n9408), .op(n7774) );
  and2_1 U9762 ( .ip1(n9425), .ip2(N4259), .op(n7773) );
  mux2_1 U9763 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[0][7] ), .s(n9391), 
        .op(n7772) );
  mux2_1 U9764 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[1][7] ), .s(n9392), 
        .op(n7771) );
  mux2_1 U9765 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[2][7] ), .s(n9393), 
        .op(n7770) );
  mux2_1 U9766 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[3][7] ), .s(n9394), 
        .op(n7769) );
  mux2_1 U9767 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[4][7] ), .s(n9395), 
        .op(n7768) );
  mux2_1 U9768 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[5][7] ), .s(n9396), 
        .op(n7767) );
  mux2_1 U9769 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[6][7] ), .s(n9397), 
        .op(n7766) );
  mux2_1 U9770 ( .ip1(addr_resp[14]), .ip2(\cache_tag_A[7][7] ), .s(n9398), 
        .op(n7765) );
  mux2_1 U9771 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[0][7] ), .s(n9399), 
        .op(n7764) );
  mux2_1 U9772 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[1][7] ), .s(n9400), 
        .op(n7763) );
  mux2_1 U9773 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[2][7] ), .s(n9401), 
        .op(n7762) );
  mux2_1 U9774 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[3][7] ), .s(n9402), 
        .op(n7761) );
  mux2_1 U9775 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[4][7] ), .s(n9403), 
        .op(n7760) );
  mux2_1 U9776 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[5][7] ), .s(n9404), 
        .op(n7759) );
  mux2_1 U9777 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[6][7] ), .s(n9405), 
        .op(n7758) );
  mux2_1 U9778 ( .ip1(addr_resp[14]), .ip2(\cache_tag_B[7][7] ), .s(n9406), 
        .op(n7757) );
  mux2_1 U9779 ( .ip1(addr_req[15]), .ip2(N4255), .s(n9408), .op(n7756) );
  and2_1 U9780 ( .ip1(n9425), .ip2(N4256), .op(n7755) );
  mux2_1 U9781 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[0][8] ), .s(n9391), 
        .op(n7754) );
  mux2_1 U9782 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[1][8] ), .s(n9392), 
        .op(n7753) );
  mux2_1 U9783 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[2][8] ), .s(n9393), 
        .op(n7752) );
  mux2_1 U9784 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[3][8] ), .s(n9394), 
        .op(n7751) );
  mux2_1 U9785 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[4][8] ), .s(n9395), 
        .op(n7750) );
  mux2_1 U9786 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[5][8] ), .s(n9396), 
        .op(n7749) );
  mux2_1 U9787 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[6][8] ), .s(n9397), 
        .op(n7748) );
  mux2_1 U9788 ( .ip1(addr_resp[15]), .ip2(\cache_tag_A[7][8] ), .s(n9398), 
        .op(n7747) );
  mux2_1 U9789 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[0][8] ), .s(n9399), 
        .op(n7746) );
  mux2_1 U9790 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[1][8] ), .s(n9400), 
        .op(n7745) );
  mux2_1 U9791 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[2][8] ), .s(n9401), 
        .op(n7744) );
  mux2_1 U9792 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[3][8] ), .s(n9402), 
        .op(n7743) );
  mux2_1 U9793 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[4][8] ), .s(n9403), 
        .op(n7742) );
  mux2_1 U9794 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[5][8] ), .s(n9404), 
        .op(n7741) );
  mux2_1 U9795 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[6][8] ), .s(n9405), 
        .op(n7740) );
  mux2_1 U9796 ( .ip1(addr_resp[15]), .ip2(\cache_tag_B[7][8] ), .s(n9406), 
        .op(n7739) );
  mux2_1 U9797 ( .ip1(addr_req[16]), .ip2(N4252), .s(n9408), .op(n7738) );
  and2_1 U9798 ( .ip1(n9425), .ip2(N4253), .op(n7737) );
  mux2_1 U9799 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[0][9] ), .s(n9391), 
        .op(n7736) );
  mux2_1 U9800 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[1][9] ), .s(n9392), 
        .op(n7735) );
  mux2_1 U9801 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[2][9] ), .s(n9393), 
        .op(n7734) );
  mux2_1 U9802 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[3][9] ), .s(n9394), 
        .op(n7733) );
  mux2_1 U9803 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[4][9] ), .s(n9395), 
        .op(n7732) );
  mux2_1 U9804 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[5][9] ), .s(n9396), 
        .op(n7731) );
  mux2_1 U9805 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[6][9] ), .s(n9397), 
        .op(n7730) );
  mux2_1 U9806 ( .ip1(addr_resp[16]), .ip2(\cache_tag_A[7][9] ), .s(n9398), 
        .op(n7729) );
  mux2_1 U9807 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[0][9] ), .s(n9399), 
        .op(n7728) );
  mux2_1 U9808 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[1][9] ), .s(n9400), 
        .op(n7727) );
  mux2_1 U9809 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[2][9] ), .s(n9401), 
        .op(n7726) );
  mux2_1 U9810 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[3][9] ), .s(n9402), 
        .op(n7725) );
  mux2_1 U9811 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[4][9] ), .s(n9403), 
        .op(n7724) );
  mux2_1 U9812 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[5][9] ), .s(n9404), 
        .op(n7723) );
  mux2_1 U9813 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[6][9] ), .s(n9405), 
        .op(n7722) );
  mux2_1 U9814 ( .ip1(addr_resp[16]), .ip2(\cache_tag_B[7][9] ), .s(n9406), 
        .op(n7721) );
  mux2_1 U9815 ( .ip1(addr_req[17]), .ip2(N4249), .s(n9408), .op(n7720) );
  and2_1 U9816 ( .ip1(n9425), .ip2(N4250), .op(n7719) );
  mux2_1 U9817 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[0][10] ), .s(n9391), 
        .op(n7718) );
  mux2_1 U9818 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[1][10] ), .s(n9392), 
        .op(n7717) );
  mux2_1 U9819 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[2][10] ), .s(n9393), 
        .op(n7716) );
  mux2_1 U9820 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[3][10] ), .s(n9394), 
        .op(n7715) );
  mux2_1 U9821 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[4][10] ), .s(n9395), 
        .op(n7714) );
  mux2_1 U9822 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[5][10] ), .s(n9396), 
        .op(n7713) );
  mux2_1 U9823 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[6][10] ), .s(n9397), 
        .op(n7712) );
  mux2_1 U9824 ( .ip1(addr_resp[17]), .ip2(\cache_tag_A[7][10] ), .s(n9398), 
        .op(n7711) );
  mux2_1 U9825 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[0][10] ), .s(n9399), 
        .op(n7710) );
  mux2_1 U9826 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[1][10] ), .s(n9400), 
        .op(n7709) );
  mux2_1 U9827 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[2][10] ), .s(n9401), 
        .op(n7708) );
  mux2_1 U9828 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[3][10] ), .s(n9402), 
        .op(n7707) );
  mux2_1 U9829 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[4][10] ), .s(n9403), 
        .op(n7706) );
  mux2_1 U9830 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[5][10] ), .s(n9404), 
        .op(n7705) );
  mux2_1 U9831 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[6][10] ), .s(n9405), 
        .op(n7704) );
  mux2_1 U9832 ( .ip1(addr_resp[17]), .ip2(\cache_tag_B[7][10] ), .s(n9406), 
        .op(n7703) );
  mux2_1 U9833 ( .ip1(addr_req[18]), .ip2(N4246), .s(n9408), .op(n7702) );
  and2_1 U9834 ( .ip1(n9425), .ip2(N4247), .op(n7701) );
  mux2_1 U9835 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[0][11] ), .s(n9391), 
        .op(n7700) );
  mux2_1 U9836 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[1][11] ), .s(n9392), 
        .op(n7699) );
  mux2_1 U9837 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[2][11] ), .s(n9393), 
        .op(n7698) );
  mux2_1 U9838 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[3][11] ), .s(n9394), 
        .op(n7697) );
  mux2_1 U9839 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[4][11] ), .s(n9395), 
        .op(n7696) );
  mux2_1 U9840 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[5][11] ), .s(n9396), 
        .op(n7695) );
  mux2_1 U9841 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[6][11] ), .s(n9397), 
        .op(n7694) );
  mux2_1 U9842 ( .ip1(addr_resp[18]), .ip2(\cache_tag_A[7][11] ), .s(n9398), 
        .op(n7693) );
  mux2_1 U9843 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[0][11] ), .s(n9399), 
        .op(n7692) );
  mux2_1 U9844 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[1][11] ), .s(n9400), 
        .op(n7691) );
  mux2_1 U9845 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[2][11] ), .s(n9401), 
        .op(n7690) );
  mux2_1 U9846 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[3][11] ), .s(n9402), 
        .op(n7689) );
  mux2_1 U9847 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[4][11] ), .s(n9403), 
        .op(n7688) );
  mux2_1 U9848 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[5][11] ), .s(n9404), 
        .op(n7687) );
  mux2_1 U9849 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[6][11] ), .s(n9405), 
        .op(n7686) );
  mux2_1 U9850 ( .ip1(addr_resp[18]), .ip2(\cache_tag_B[7][11] ), .s(n9406), 
        .op(n7685) );
  mux2_1 U9851 ( .ip1(addr_req[19]), .ip2(N4243), .s(n9408), .op(n7684) );
  and2_1 U9852 ( .ip1(n9425), .ip2(N4244), .op(n7683) );
  mux2_1 U9853 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[0][12] ), .s(n9391), 
        .op(n7682) );
  mux2_1 U9854 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[1][12] ), .s(n9392), 
        .op(n7681) );
  mux2_1 U9855 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[2][12] ), .s(n9393), 
        .op(n7680) );
  mux2_1 U9856 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[3][12] ), .s(n9394), 
        .op(n7679) );
  mux2_1 U9857 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[4][12] ), .s(n9395), 
        .op(n7678) );
  mux2_1 U9858 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[5][12] ), .s(n9396), 
        .op(n7677) );
  mux2_1 U9859 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[6][12] ), .s(n9397), 
        .op(n7676) );
  mux2_1 U9860 ( .ip1(addr_resp[19]), .ip2(\cache_tag_A[7][12] ), .s(n9398), 
        .op(n7675) );
  mux2_1 U9861 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[0][12] ), .s(n9399), 
        .op(n7674) );
  mux2_1 U9862 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[1][12] ), .s(n9400), 
        .op(n7673) );
  mux2_1 U9863 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[2][12] ), .s(n9401), 
        .op(n7672) );
  mux2_1 U9864 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[3][12] ), .s(n9402), 
        .op(n7671) );
  mux2_1 U9865 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[4][12] ), .s(n9403), 
        .op(n7670) );
  mux2_1 U9866 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[5][12] ), .s(n9404), 
        .op(n7669) );
  mux2_1 U9867 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[6][12] ), .s(n9405), 
        .op(n7668) );
  mux2_1 U9868 ( .ip1(addr_resp[19]), .ip2(\cache_tag_B[7][12] ), .s(n9406), 
        .op(n7667) );
  mux2_1 U9869 ( .ip1(addr_req[20]), .ip2(N4240), .s(n9408), .op(n7666) );
  and2_1 U9870 ( .ip1(n9425), .ip2(N4241), .op(n7665) );
  mux2_1 U9871 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[0][13] ), .s(n9391), 
        .op(n7664) );
  mux2_1 U9872 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[1][13] ), .s(n9392), 
        .op(n7663) );
  mux2_1 U9873 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[2][13] ), .s(n9393), 
        .op(n7662) );
  mux2_1 U9874 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[3][13] ), .s(n9394), 
        .op(n7661) );
  mux2_1 U9875 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[4][13] ), .s(n9395), 
        .op(n7660) );
  mux2_1 U9876 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[5][13] ), .s(n9396), 
        .op(n7659) );
  mux2_1 U9877 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[6][13] ), .s(n9397), 
        .op(n7658) );
  mux2_1 U9878 ( .ip1(addr_resp[20]), .ip2(\cache_tag_A[7][13] ), .s(n9398), 
        .op(n7657) );
  mux2_1 U9879 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[0][13] ), .s(n9399), 
        .op(n7656) );
  mux2_1 U9880 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[1][13] ), .s(n9400), 
        .op(n7655) );
  mux2_1 U9881 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[2][13] ), .s(n9401), 
        .op(n7654) );
  mux2_1 U9882 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[3][13] ), .s(n9402), 
        .op(n7653) );
  mux2_1 U9883 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[4][13] ), .s(n9403), 
        .op(n7652) );
  mux2_1 U9884 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[5][13] ), .s(n9404), 
        .op(n7651) );
  mux2_1 U9885 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[6][13] ), .s(n9405), 
        .op(n7650) );
  mux2_1 U9886 ( .ip1(addr_resp[20]), .ip2(\cache_tag_B[7][13] ), .s(n9406), 
        .op(n7649) );
  mux2_1 U9887 ( .ip1(addr_req[21]), .ip2(N4237), .s(n9425), .op(n7648) );
  and2_1 U9888 ( .ip1(n9408), .ip2(N4238), .op(n7647) );
  mux2_1 U9889 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[0][14] ), .s(n9391), 
        .op(n7646) );
  mux2_1 U9890 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[1][14] ), .s(n9392), 
        .op(n7645) );
  mux2_1 U9891 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[2][14] ), .s(n9393), 
        .op(n7644) );
  mux2_1 U9892 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[3][14] ), .s(n9394), 
        .op(n7643) );
  mux2_1 U9893 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[4][14] ), .s(n9395), 
        .op(n7642) );
  mux2_1 U9894 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[5][14] ), .s(n9396), 
        .op(n7641) );
  mux2_1 U9895 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[6][14] ), .s(n9397), 
        .op(n7640) );
  mux2_1 U9896 ( .ip1(addr_resp[21]), .ip2(\cache_tag_A[7][14] ), .s(n9398), 
        .op(n7639) );
  mux2_1 U9897 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[0][14] ), .s(n9399), 
        .op(n7638) );
  mux2_1 U9898 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[1][14] ), .s(n9400), 
        .op(n7637) );
  mux2_1 U9899 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[2][14] ), .s(n9401), 
        .op(n7636) );
  mux2_1 U9900 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[3][14] ), .s(n9402), 
        .op(n7635) );
  mux2_1 U9901 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[4][14] ), .s(n9403), 
        .op(n7634) );
  mux2_1 U9902 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[5][14] ), .s(n9404), 
        .op(n7633) );
  mux2_1 U9903 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[6][14] ), .s(n9405), 
        .op(n7632) );
  mux2_1 U9904 ( .ip1(addr_resp[21]), .ip2(\cache_tag_B[7][14] ), .s(n9406), 
        .op(n7631) );
  mux2_1 U9905 ( .ip1(addr_req[22]), .ip2(N4234), .s(n9408), .op(n7630) );
  and2_1 U9906 ( .ip1(n9408), .ip2(N4235), .op(n7629) );
  mux2_1 U9907 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[0][15] ), .s(n9391), 
        .op(n7628) );
  mux2_1 U9908 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[1][15] ), .s(n9392), 
        .op(n7627) );
  mux2_1 U9909 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[2][15] ), .s(n9393), 
        .op(n7626) );
  mux2_1 U9910 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[3][15] ), .s(n9394), 
        .op(n7625) );
  mux2_1 U9911 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[4][15] ), .s(n9395), 
        .op(n7624) );
  mux2_1 U9912 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[5][15] ), .s(n9396), 
        .op(n7623) );
  mux2_1 U9913 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[6][15] ), .s(n9397), 
        .op(n7622) );
  mux2_1 U9914 ( .ip1(addr_resp[22]), .ip2(\cache_tag_A[7][15] ), .s(n9398), 
        .op(n7621) );
  mux2_1 U9915 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[0][15] ), .s(n9399), 
        .op(n7620) );
  mux2_1 U9916 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[1][15] ), .s(n9400), 
        .op(n7619) );
  mux2_1 U9917 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[2][15] ), .s(n9401), 
        .op(n7618) );
  mux2_1 U9918 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[3][15] ), .s(n9402), 
        .op(n7617) );
  mux2_1 U9919 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[4][15] ), .s(n9403), 
        .op(n7616) );
  mux2_1 U9920 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[5][15] ), .s(n9404), 
        .op(n7615) );
  mux2_1 U9921 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[6][15] ), .s(n9405), 
        .op(n7614) );
  mux2_1 U9922 ( .ip1(addr_resp[22]), .ip2(\cache_tag_B[7][15] ), .s(n9406), 
        .op(n7613) );
  mux2_1 U9923 ( .ip1(addr_req[23]), .ip2(N4231), .s(n9408), .op(n7612) );
  and2_1 U9924 ( .ip1(n9408), .ip2(N4232), .op(n7611) );
  mux2_1 U9925 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[0][16] ), .s(n9409), 
        .op(n7610) );
  mux2_1 U9926 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[1][16] ), .s(n9410), 
        .op(n7609) );
  mux2_1 U9927 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[2][16] ), .s(n9411), 
        .op(n7608) );
  mux2_1 U9928 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[3][16] ), .s(n9412), 
        .op(n7607) );
  mux2_1 U9929 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[4][16] ), .s(n9413), 
        .op(n7606) );
  mux2_1 U9930 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[5][16] ), .s(n9414), 
        .op(n7605) );
  mux2_1 U9931 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[6][16] ), .s(n9415), 
        .op(n7604) );
  mux2_1 U9932 ( .ip1(addr_resp[23]), .ip2(\cache_tag_A[7][16] ), .s(n9416), 
        .op(n7603) );
  mux2_1 U9933 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[0][16] ), .s(n9417), 
        .op(n7602) );
  mux2_1 U9934 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[1][16] ), .s(n9418), 
        .op(n7601) );
  mux2_1 U9935 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[2][16] ), .s(n9419), 
        .op(n7600) );
  mux2_1 U9936 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[3][16] ), .s(n9420), 
        .op(n7599) );
  mux2_1 U9937 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[4][16] ), .s(n9421), 
        .op(n7598) );
  mux2_1 U9938 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[5][16] ), .s(n9422), 
        .op(n7597) );
  mux2_1 U9939 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[6][16] ), .s(n9423), 
        .op(n7596) );
  mux2_1 U9940 ( .ip1(addr_resp[23]), .ip2(\cache_tag_B[7][16] ), .s(n9424), 
        .op(n7595) );
  mux2_1 U9941 ( .ip1(addr_req[24]), .ip2(N4228), .s(n9408), .op(n7594) );
  and2_1 U9942 ( .ip1(n9408), .ip2(N4229), .op(n7593) );
  mux2_1 U9943 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[0][17] ), .s(n9391), 
        .op(n7592) );
  mux2_1 U9944 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[1][17] ), .s(n9392), 
        .op(n7591) );
  mux2_1 U9945 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[2][17] ), .s(n9393), 
        .op(n7590) );
  mux2_1 U9946 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[3][17] ), .s(n9394), 
        .op(n7589) );
  mux2_1 U9947 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[4][17] ), .s(n9395), 
        .op(n7588) );
  mux2_1 U9948 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[5][17] ), .s(n9396), 
        .op(n7587) );
  mux2_1 U9949 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[6][17] ), .s(n9397), 
        .op(n7586) );
  mux2_1 U9950 ( .ip1(addr_resp[24]), .ip2(\cache_tag_A[7][17] ), .s(n9398), 
        .op(n7585) );
  mux2_1 U9951 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[0][17] ), .s(n9399), 
        .op(n7584) );
  mux2_1 U9952 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[1][17] ), .s(n9400), 
        .op(n7583) );
  mux2_1 U9953 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[2][17] ), .s(n9401), 
        .op(n7582) );
  mux2_1 U9954 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[3][17] ), .s(n9402), 
        .op(n7581) );
  mux2_1 U9955 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[4][17] ), .s(n9403), 
        .op(n7580) );
  mux2_1 U9956 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[5][17] ), .s(n9404), 
        .op(n7579) );
  mux2_1 U9957 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[6][17] ), .s(n9405), 
        .op(n7578) );
  mux2_1 U9958 ( .ip1(addr_resp[24]), .ip2(\cache_tag_B[7][17] ), .s(n9406), 
        .op(n7577) );
  mux2_1 U9959 ( .ip1(addr_req[25]), .ip2(N4225), .s(n9425), .op(n7576) );
  and2_1 U9960 ( .ip1(n9408), .ip2(N4226), .op(n7575) );
  mux2_1 U9961 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[0][18] ), .s(n9409), 
        .op(n7574) );
  mux2_1 U9962 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[1][18] ), .s(n9410), 
        .op(n7573) );
  mux2_1 U9963 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[2][18] ), .s(n9411), 
        .op(n7572) );
  mux2_1 U9964 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[3][18] ), .s(n9412), 
        .op(n7571) );
  mux2_1 U9965 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[4][18] ), .s(n9413), 
        .op(n7570) );
  mux2_1 U9966 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[5][18] ), .s(n9414), 
        .op(n7569) );
  mux2_1 U9967 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[6][18] ), .s(n9415), 
        .op(n7568) );
  mux2_1 U9968 ( .ip1(addr_resp[25]), .ip2(\cache_tag_A[7][18] ), .s(n9416), 
        .op(n7567) );
  mux2_1 U9969 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[0][18] ), .s(n9417), 
        .op(n7566) );
  mux2_1 U9970 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[1][18] ), .s(n9418), 
        .op(n7565) );
  mux2_1 U9971 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[2][18] ), .s(n9419), 
        .op(n7564) );
  mux2_1 U9972 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[3][18] ), .s(n9420), 
        .op(n7563) );
  mux2_1 U9973 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[4][18] ), .s(n9421), 
        .op(n7562) );
  mux2_1 U9974 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[5][18] ), .s(n9422), 
        .op(n7561) );
  mux2_1 U9975 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[6][18] ), .s(n9423), 
        .op(n7560) );
  mux2_1 U9976 ( .ip1(addr_resp[25]), .ip2(\cache_tag_B[7][18] ), .s(n9424), 
        .op(n7559) );
  mux2_1 U9977 ( .ip1(addr_req[26]), .ip2(N4222), .s(n9408), .op(n7558) );
  and2_1 U9978 ( .ip1(n9408), .ip2(N4223), .op(n7557) );
  mux2_1 U9979 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[0][19] ), .s(n9391), 
        .op(n7556) );
  mux2_1 U9980 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[1][19] ), .s(n9392), 
        .op(n7555) );
  mux2_1 U9981 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[2][19] ), .s(n9393), 
        .op(n7554) );
  mux2_1 U9982 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[3][19] ), .s(n9394), 
        .op(n7553) );
  mux2_1 U9983 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[4][19] ), .s(n9395), 
        .op(n7552) );
  mux2_1 U9984 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[5][19] ), .s(n9396), 
        .op(n7551) );
  mux2_1 U9985 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[6][19] ), .s(n9397), 
        .op(n7550) );
  mux2_1 U9986 ( .ip1(addr_resp[26]), .ip2(\cache_tag_A[7][19] ), .s(n9398), 
        .op(n7549) );
  mux2_1 U9987 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[0][19] ), .s(n9399), 
        .op(n7548) );
  mux2_1 U9988 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[1][19] ), .s(n9400), 
        .op(n7547) );
  mux2_1 U9989 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[2][19] ), .s(n9401), 
        .op(n7546) );
  mux2_1 U9990 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[3][19] ), .s(n9402), 
        .op(n7545) );
  mux2_1 U9991 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[4][19] ), .s(n9403), 
        .op(n7544) );
  mux2_1 U9992 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[5][19] ), .s(n9404), 
        .op(n7543) );
  mux2_1 U9993 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[6][19] ), .s(n9405), 
        .op(n7542) );
  mux2_1 U9994 ( .ip1(addr_resp[26]), .ip2(\cache_tag_B[7][19] ), .s(n9406), 
        .op(n7541) );
  mux2_1 U9995 ( .ip1(addr_req[27]), .ip2(N4219), .s(n9407), .op(n7540) );
  and2_1 U9996 ( .ip1(n9408), .ip2(N4220), .op(n7539) );
  mux2_1 U9997 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[0][20] ), .s(n9409), 
        .op(n7538) );
  mux2_1 U9998 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[1][20] ), .s(n9410), 
        .op(n7537) );
  mux2_1 U9999 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[2][20] ), .s(n9411), 
        .op(n7536) );
  mux2_1 U10000 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[3][20] ), .s(n9412), 
        .op(n7535) );
  mux2_1 U10001 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[4][20] ), .s(n9413), 
        .op(n7534) );
  mux2_1 U10002 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[5][20] ), .s(n9414), 
        .op(n7533) );
  mux2_1 U10003 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[6][20] ), .s(n9415), 
        .op(n7532) );
  mux2_1 U10004 ( .ip1(addr_resp[27]), .ip2(\cache_tag_A[7][20] ), .s(n9416), 
        .op(n7531) );
  mux2_1 U10005 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[0][20] ), .s(n9417), 
        .op(n7530) );
  mux2_1 U10006 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[1][20] ), .s(n9418), 
        .op(n7529) );
  mux2_1 U10007 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[2][20] ), .s(n9419), 
        .op(n7528) );
  mux2_1 U10008 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[3][20] ), .s(n9420), 
        .op(n7527) );
  mux2_1 U10009 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[4][20] ), .s(n9421), 
        .op(n7526) );
  mux2_1 U10010 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[5][20] ), .s(n9422), 
        .op(n7525) );
  mux2_1 U10011 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[6][20] ), .s(n9423), 
        .op(n7524) );
  mux2_1 U10012 ( .ip1(addr_resp[27]), .ip2(\cache_tag_B[7][20] ), .s(n9424), 
        .op(n7523) );
  mux2_1 U10013 ( .ip1(addr_req[28]), .ip2(N4216), .s(n9425), .op(n7522) );
  and2_1 U10014 ( .ip1(n9408), .ip2(N4217), .op(n7521) );
  mux2_1 U10015 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[0][21] ), .s(n9391), 
        .op(n7520) );
  mux2_1 U10016 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[1][21] ), .s(n9392), 
        .op(n7519) );
  mux2_1 U10017 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[2][21] ), .s(n9393), 
        .op(n7518) );
  mux2_1 U10018 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[3][21] ), .s(n9394), 
        .op(n7517) );
  mux2_1 U10019 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[4][21] ), .s(n9395), 
        .op(n7516) );
  mux2_1 U10020 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[5][21] ), .s(n9396), 
        .op(n7515) );
  mux2_1 U10021 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[6][21] ), .s(n9397), 
        .op(n7514) );
  mux2_1 U10022 ( .ip1(addr_resp[28]), .ip2(\cache_tag_A[7][21] ), .s(n9398), 
        .op(n7513) );
  mux2_1 U10023 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[0][21] ), .s(n9399), 
        .op(n7512) );
  mux2_1 U10024 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[1][21] ), .s(n9400), 
        .op(n7511) );
  mux2_1 U10025 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[2][21] ), .s(n9401), 
        .op(n7510) );
  mux2_1 U10026 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[3][21] ), .s(n9402), 
        .op(n7509) );
  mux2_1 U10027 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[4][21] ), .s(n9403), 
        .op(n7508) );
  mux2_1 U10028 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[5][21] ), .s(n9404), 
        .op(n7507) );
  mux2_1 U10029 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[6][21] ), .s(n9405), 
        .op(n7506) );
  mux2_1 U10030 ( .ip1(addr_resp[28]), .ip2(\cache_tag_B[7][21] ), .s(n9406), 
        .op(n7505) );
  mux2_1 U10031 ( .ip1(addr_req[29]), .ip2(N4213), .s(n9407), .op(n7504) );
  and2_1 U10032 ( .ip1(n9408), .ip2(N4214), .op(n7503) );
  mux2_1 U10033 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[0][22] ), .s(n9409), 
        .op(n7502) );
  mux2_1 U10034 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[1][22] ), .s(n9410), 
        .op(n7501) );
  mux2_1 U10035 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[2][22] ), .s(n9411), 
        .op(n7500) );
  mux2_1 U10036 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[3][22] ), .s(n9412), 
        .op(n7499) );
  mux2_1 U10037 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[4][22] ), .s(n9413), 
        .op(n7498) );
  mux2_1 U10038 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[5][22] ), .s(n9414), 
        .op(n7497) );
  mux2_1 U10039 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[6][22] ), .s(n9415), 
        .op(n7496) );
  mux2_1 U10040 ( .ip1(addr_resp[29]), .ip2(\cache_tag_A[7][22] ), .s(n9416), 
        .op(n7495) );
  mux2_1 U10041 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[0][22] ), .s(n9417), 
        .op(n7494) );
  mux2_1 U10042 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[1][22] ), .s(n9418), 
        .op(n7493) );
  mux2_1 U10043 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[2][22] ), .s(n9419), 
        .op(n7492) );
  mux2_1 U10044 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[3][22] ), .s(n9420), 
        .op(n7491) );
  mux2_1 U10045 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[4][22] ), .s(n9421), 
        .op(n7490) );
  mux2_1 U10046 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[5][22] ), .s(n9422), 
        .op(n7489) );
  mux2_1 U10047 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[6][22] ), .s(n9423), 
        .op(n7488) );
  mux2_1 U10048 ( .ip1(addr_resp[29]), .ip2(\cache_tag_B[7][22] ), .s(n9424), 
        .op(n7487) );
  mux2_1 U10049 ( .ip1(addr_req[30]), .ip2(N4210), .s(n9407), .op(n7486) );
  and2_1 U10050 ( .ip1(n9408), .ip2(N4211), .op(n7485) );
  mux2_1 U10051 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[0][23] ), .s(n9391), 
        .op(n7484) );
  mux2_1 U10052 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[1][23] ), .s(n9392), 
        .op(n7483) );
  mux2_1 U10053 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[2][23] ), .s(n9393), 
        .op(n7482) );
  mux2_1 U10054 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[3][23] ), .s(n9394), 
        .op(n7481) );
  mux2_1 U10055 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[4][23] ), .s(n9395), 
        .op(n7480) );
  mux2_1 U10056 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[5][23] ), .s(n9396), 
        .op(n7479) );
  mux2_1 U10057 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[6][23] ), .s(n9397), 
        .op(n7478) );
  mux2_1 U10058 ( .ip1(addr_resp[30]), .ip2(\cache_tag_A[7][23] ), .s(n9398), 
        .op(n7477) );
  mux2_1 U10059 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[0][23] ), .s(n9399), 
        .op(n7476) );
  mux2_1 U10060 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[1][23] ), .s(n9400), 
        .op(n7475) );
  mux2_1 U10061 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[2][23] ), .s(n9401), 
        .op(n7474) );
  mux2_1 U10062 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[3][23] ), .s(n9402), 
        .op(n7473) );
  mux2_1 U10063 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[4][23] ), .s(n9403), 
        .op(n7472) );
  mux2_1 U10064 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[5][23] ), .s(n9404), 
        .op(n7471) );
  mux2_1 U10065 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[6][23] ), .s(n9405), 
        .op(n7470) );
  mux2_1 U10066 ( .ip1(addr_resp[30]), .ip2(\cache_tag_B[7][23] ), .s(n9406), 
        .op(n7469) );
  mux2_1 U10067 ( .ip1(addr_req[31]), .ip2(N4207), .s(n9407), .op(n7468) );
  and2_1 U10068 ( .ip1(n9408), .ip2(N4208), .op(n7467) );
  mux2_1 U10069 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[0][24] ), .s(n9409), 
        .op(n7466) );
  mux2_1 U10070 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[1][24] ), .s(n9410), 
        .op(n7465) );
  mux2_1 U10071 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[2][24] ), .s(n9411), 
        .op(n7464) );
  mux2_1 U10072 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[3][24] ), .s(n9412), 
        .op(n7463) );
  mux2_1 U10073 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[4][24] ), .s(n9413), 
        .op(n7462) );
  mux2_1 U10074 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[5][24] ), .s(n9414), 
        .op(n7461) );
  mux2_1 U10075 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[6][24] ), .s(n9415), 
        .op(n7460) );
  mux2_1 U10076 ( .ip1(addr_resp[31]), .ip2(\cache_tag_A[7][24] ), .s(n9416), 
        .op(n7459) );
  mux2_1 U10077 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[0][24] ), .s(n9417), 
        .op(n7458) );
  mux2_1 U10078 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[1][24] ), .s(n9418), 
        .op(n7457) );
  mux2_1 U10079 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[2][24] ), .s(n9419), 
        .op(n7456) );
  mux2_1 U10080 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[3][24] ), .s(n9420), 
        .op(n7455) );
  mux2_1 U10081 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[4][24] ), .s(n9421), 
        .op(n7454) );
  mux2_1 U10082 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[5][24] ), .s(n9422), 
        .op(n7453) );
  mux2_1 U10083 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[6][24] ), .s(n9423), 
        .op(n7452) );
  mux2_1 U10084 ( .ip1(addr_resp[31]), .ip2(\cache_tag_B[7][24] ), .s(n9424), 
        .op(n7451) );
  nor2_1 U10085 ( .ip1(n12618), .ip2(n9425), .op(n9426) );
  buf_1 U10086 ( .ip(n9426), .op(n9427) );
  mux2_1 U10087 ( .ip1(iCache_data_wr[0]), .ip2(data_wr[0]), .s(n9427), .op(
        n7450) );
  mux2_1 U10088 ( .ip1(iCache_data_wr[1]), .ip2(data_wr[1]), .s(n9426), .op(
        n7449) );
  mux2_1 U10089 ( .ip1(iCache_data_wr[2]), .ip2(data_wr[2]), .s(n9426), .op(
        n7448) );
  mux2_1 U10090 ( .ip1(iCache_data_wr[3]), .ip2(data_wr[3]), .s(n9426), .op(
        n7447) );
  mux2_1 U10091 ( .ip1(iCache_data_wr[4]), .ip2(data_wr[4]), .s(n9426), .op(
        n7446) );
  mux2_1 U10092 ( .ip1(iCache_data_wr[5]), .ip2(data_wr[5]), .s(n9426), .op(
        n7445) );
  mux2_1 U10093 ( .ip1(iCache_data_wr[6]), .ip2(data_wr[6]), .s(n9426), .op(
        n7444) );
  mux2_1 U10094 ( .ip1(iCache_data_wr[7]), .ip2(data_wr[7]), .s(n9426), .op(
        n7443) );
  mux2_1 U10095 ( .ip1(iCache_data_wr[8]), .ip2(data_wr[8]), .s(n9426), .op(
        n7442) );
  mux2_1 U10096 ( .ip1(iCache_data_wr[9]), .ip2(data_wr[9]), .s(n9427), .op(
        n7441) );
  mux2_1 U10097 ( .ip1(iCache_data_wr[10]), .ip2(data_wr[10]), .s(n9427), .op(
        n7440) );
  mux2_1 U10098 ( .ip1(iCache_data_wr[11]), .ip2(data_wr[11]), .s(n9426), .op(
        n7439) );
  mux2_1 U10099 ( .ip1(iCache_data_wr[12]), .ip2(data_wr[12]), .s(n9426), .op(
        n7438) );
  mux2_1 U10100 ( .ip1(iCache_data_wr[13]), .ip2(data_wr[13]), .s(n9426), .op(
        n7437) );
  mux2_1 U10101 ( .ip1(iCache_data_wr[14]), .ip2(data_wr[14]), .s(n9426), .op(
        n7436) );
  mux2_1 U10102 ( .ip1(iCache_data_wr[15]), .ip2(data_wr[15]), .s(n9426), .op(
        n7435) );
  mux2_1 U10103 ( .ip1(iCache_data_wr[16]), .ip2(data_wr[16]), .s(n9426), .op(
        n7434) );
  mux2_1 U10104 ( .ip1(iCache_data_wr[17]), .ip2(data_wr[17]), .s(n9426), .op(
        n7433) );
  mux2_1 U10105 ( .ip1(iCache_data_wr[18]), .ip2(data_wr[18]), .s(n9426), .op(
        n7432) );
  mux2_1 U10106 ( .ip1(iCache_data_wr[19]), .ip2(data_wr[19]), .s(n9426), .op(
        n7431) );
  mux2_1 U10107 ( .ip1(iCache_data_wr[20]), .ip2(data_wr[20]), .s(n9426), .op(
        n7430) );
  mux2_1 U10108 ( .ip1(iCache_data_wr[21]), .ip2(data_wr[21]), .s(n9426), .op(
        n7429) );
  mux2_1 U10109 ( .ip1(iCache_data_wr[22]), .ip2(data_wr[22]), .s(n9426), .op(
        n7428) );
  mux2_1 U10110 ( .ip1(iCache_data_wr[23]), .ip2(data_wr[23]), .s(n9426), .op(
        n7427) );
  mux2_1 U10111 ( .ip1(iCache_data_wr[24]), .ip2(data_wr[24]), .s(n9427), .op(
        n7426) );
  mux2_1 U10112 ( .ip1(iCache_data_wr[25]), .ip2(data_wr[25]), .s(n9427), .op(
        n7425) );
  mux2_1 U10113 ( .ip1(iCache_data_wr[26]), .ip2(data_wr[26]), .s(n9427), .op(
        n7424) );
  mux2_1 U10114 ( .ip1(iCache_data_wr[27]), .ip2(data_wr[27]), .s(n9427), .op(
        n7423) );
  mux2_1 U10115 ( .ip1(iCache_data_wr[28]), .ip2(data_wr[28]), .s(n9427), .op(
        n7422) );
  mux2_1 U10116 ( .ip1(iCache_data_wr[29]), .ip2(data_wr[29]), .s(n9427), .op(
        n7421) );
  mux2_1 U10117 ( .ip1(iCache_data_wr[30]), .ip2(data_wr[30]), .s(n9427), .op(
        n7420) );
  mux2_1 U10118 ( .ip1(iCache_data_wr[31]), .ip2(data_wr[31]), .s(n9427), .op(
        n7419) );
  buf_1 U10119 ( .ip(n13294), .op(n9872) );
  and2_1 U10120 ( .ip1(n9872), .ip2(rd_temp), .op(n10378) );
  inv_1 U10121 ( .ip(N4205), .op(n9428) );
  nor2_1 U10122 ( .ip1(n10378), .ip2(n9428), .op(n7418) );
  inv_1 U10123 ( .ip(N4202), .op(n9429) );
  nor2_1 U10124 ( .ip1(n10378), .ip2(n9429), .op(n7417) );
  inv_1 U10125 ( .ip(N4199), .op(n9430) );
  nor2_1 U10126 ( .ip1(n10378), .ip2(n9430), .op(n7416) );
  buf_1 U10127 ( .ip(n10378), .op(n11472) );
  inv_1 U10128 ( .ip(N4196), .op(n9431) );
  nor2_1 U10129 ( .ip1(n11472), .ip2(n9431), .op(n7415) );
  buf_1 U10130 ( .ip(n10378), .op(n12599) );
  inv_1 U10131 ( .ip(N4193), .op(n9432) );
  nor2_1 U10132 ( .ip1(n12599), .ip2(n9432), .op(n7414) );
  inv_1 U10133 ( .ip(N4190), .op(n9433) );
  nor2_1 U10134 ( .ip1(n10378), .ip2(n9433), .op(n7413) );
  inv_1 U10135 ( .ip(N4187), .op(n9434) );
  nor2_1 U10136 ( .ip1(n11472), .ip2(n9434), .op(n7412) );
  inv_1 U10137 ( .ip(N4184), .op(n9435) );
  nor2_1 U10138 ( .ip1(n12599), .ip2(n9435), .op(n7411) );
  inv_1 U10139 ( .ip(N4181), .op(n9436) );
  nor2_1 U10140 ( .ip1(n10378), .ip2(n9436), .op(n7410) );
  inv_1 U10141 ( .ip(N4178), .op(n9437) );
  nor2_1 U10142 ( .ip1(n11472), .ip2(n9437), .op(n7409) );
  inv_1 U10143 ( .ip(N4175), .op(n9438) );
  nor2_1 U10144 ( .ip1(n12599), .ip2(n9438), .op(n7408) );
  inv_1 U10145 ( .ip(N4172), .op(n9439) );
  nor2_1 U10146 ( .ip1(n10378), .ip2(n9439), .op(n7407) );
  inv_1 U10147 ( .ip(N4169), .op(n9440) );
  nor2_1 U10148 ( .ip1(n11472), .ip2(n9440), .op(n7406) );
  inv_1 U10149 ( .ip(N4166), .op(n9441) );
  nor2_1 U10150 ( .ip1(n12599), .ip2(n9441), .op(n7405) );
  inv_1 U10151 ( .ip(N4163), .op(n9442) );
  nor2_1 U10152 ( .ip1(n10378), .ip2(n9442), .op(n7404) );
  inv_1 U10153 ( .ip(N4160), .op(n9443) );
  nor2_1 U10154 ( .ip1(n10378), .ip2(n9443), .op(n7403) );
  inv_1 U10155 ( .ip(N4157), .op(n9444) );
  nor2_1 U10156 ( .ip1(n10378), .ip2(n9444), .op(n7402) );
  inv_1 U10157 ( .ip(N4154), .op(n9445) );
  nor2_1 U10158 ( .ip1(n10378), .ip2(n9445), .op(n7401) );
  inv_1 U10159 ( .ip(N4151), .op(n9446) );
  nor2_1 U10160 ( .ip1(n10378), .ip2(n9446), .op(n7400) );
  inv_1 U10161 ( .ip(N4148), .op(n9447) );
  nor2_1 U10162 ( .ip1(n10378), .ip2(n9447), .op(n7399) );
  inv_1 U10163 ( .ip(N4145), .op(n9448) );
  nor2_1 U10164 ( .ip1(n10378), .ip2(n9448), .op(n7398) );
  inv_1 U10165 ( .ip(N4142), .op(n9449) );
  nor2_1 U10166 ( .ip1(n10378), .ip2(n9449), .op(n7397) );
  inv_1 U10167 ( .ip(N4139), .op(n9450) );
  nor2_1 U10168 ( .ip1(n10378), .ip2(n9450), .op(n7396) );
  inv_1 U10169 ( .ip(N4136), .op(n9451) );
  nor2_1 U10170 ( .ip1(n10378), .ip2(n9451), .op(n7395) );
  inv_1 U10171 ( .ip(N4133), .op(n9452) );
  nor2_1 U10172 ( .ip1(n10378), .ip2(n9452), .op(n7394) );
  inv_1 U10173 ( .ip(N4130), .op(n9453) );
  nor2_1 U10174 ( .ip1(n10378), .ip2(n9453), .op(n7393) );
  inv_1 U10175 ( .ip(N4127), .op(n9454) );
  nor2_1 U10176 ( .ip1(n10378), .ip2(n9454), .op(n7392) );
  inv_1 U10177 ( .ip(N4124), .op(n9455) );
  nor2_1 U10178 ( .ip1(n10378), .ip2(n9455), .op(n7391) );
  inv_1 U10179 ( .ip(N4121), .op(n9456) );
  nor2_1 U10180 ( .ip1(n10378), .ip2(n9456), .op(n7390) );
  inv_1 U10181 ( .ip(N4118), .op(n9457) );
  nor2_1 U10182 ( .ip1(n10378), .ip2(n9457), .op(n7389) );
  inv_1 U10183 ( .ip(N4115), .op(n9458) );
  nor2_1 U10184 ( .ip1(n10378), .ip2(n9458), .op(n7388) );
  inv_1 U10185 ( .ip(N4112), .op(n9459) );
  nor2_1 U10186 ( .ip1(n10378), .ip2(n9459), .op(n7387) );
  nand2_1 U10187 ( .ip1(n13191), .ip2(n13189), .op(n13200) );
  nand2_1 U10188 ( .ip1(mem_data_cnt[2]), .ip2(n13200), .op(n13193) );
  mux2_1 U10189 ( .ip1(n9701), .ip2(mem_data_cnt[3]), .s(n13193), .op(n7386)
         );
  mux2_1 U10190 ( .ip1(mem_data_cnt[2]), .ip2(n9700), .s(n13200), .op(n7385)
         );
  nand2_1 U10191 ( .ip1(data_rd_mem[25]), .ip2(n13295), .op(n9461) );
  nand2_1 U10192 ( .ip1(iCache_data_wr[25]), .ip2(n9872), .op(n9460) );
  nand2_1 U10193 ( .ip1(n9461), .ip2(n9460), .op(n9838) );
  nor3_1 U10194 ( .ip1(SelectWay), .ip2(mem_data_cnt[3]), .ip3(mem_data_cnt[2]), .op(n13180) );
  nand2_1 U10195 ( .ip1(n13180), .ip2(n9619), .op(n9546) );
  inv_1 U10196 ( .ip(addr_resp[3]), .op(n9704) );
  inv_1 U10197 ( .ip(addr_resp[2]), .op(n9705) );
  nand2_1 U10198 ( .ip1(n9704), .ip2(n9705), .op(n9924) );
  inv_1 U10199 ( .ip(n9924), .op(n9687) );
  inv_1 U10200 ( .ip(addr_resp[28]), .op(n9463) );
  mux2_1 U10201 ( .ip1(addr_resp[28]), .ip2(n9463), .s(n9462), .op(n9473) );
  inv_1 U10202 ( .ip(addr_resp[21]), .op(n9465) );
  mux2_1 U10203 ( .ip1(addr_resp[21]), .ip2(n9465), .s(n9464), .op(n9472) );
  inv_1 U10204 ( .ip(addr_resp[15]), .op(n9467) );
  mux2_1 U10205 ( .ip1(addr_resp[15]), .ip2(n9467), .s(n9466), .op(n9471) );
  inv_1 U10206 ( .ip(addr_resp[24]), .op(n9469) );
  mux2_1 U10207 ( .ip1(addr_resp[24]), .ip2(n9469), .s(n9468), .op(n9470) );
  nor4_1 U10208 ( .ip1(n9473), .ip2(n9472), .ip3(n9471), .ip4(n9470), .op(
        n9543) );
  inv_1 U10209 ( .ip(addr_resp[25]), .op(n9475) );
  mux2_1 U10210 ( .ip1(n9475), .ip2(addr_resp[25]), .s(n9474), .op(n9542) );
  inv_1 U10211 ( .ip(addr_resp[30]), .op(n9477) );
  mux2_1 U10212 ( .ip1(addr_resp[30]), .ip2(n9477), .s(n9476), .op(n9487) );
  inv_1 U10213 ( .ip(addr_resp[19]), .op(n9479) );
  mux2_1 U10214 ( .ip1(addr_resp[19]), .ip2(n9479), .s(n9478), .op(n9486) );
  inv_1 U10215 ( .ip(addr_resp[26]), .op(n9481) );
  mux2_1 U10216 ( .ip1(addr_resp[26]), .ip2(n9481), .s(n9480), .op(n9485) );
  inv_1 U10217 ( .ip(addr_resp[14]), .op(n9483) );
  mux2_1 U10218 ( .ip1(addr_resp[14]), .ip2(n9483), .s(n9482), .op(n9484) );
  nor4_1 U10219 ( .ip1(n9487), .ip2(n9486), .ip3(n9485), .ip4(n9484), .op(
        n9541) );
  inv_1 U10220 ( .ip(addr_resp[18]), .op(n9489) );
  mux2_1 U10221 ( .ip1(n9489), .ip2(addr_resp[18]), .s(n9488), .op(n9499) );
  inv_1 U10222 ( .ip(addr_resp[12]), .op(n9491) );
  mux2_1 U10223 ( .ip1(n9491), .ip2(addr_resp[12]), .s(n9490), .op(n9498) );
  inv_1 U10224 ( .ip(addr_resp[8]), .op(n9493) );
  mux2_1 U10225 ( .ip1(n9493), .ip2(addr_resp[8]), .s(n9492), .op(n9497) );
  inv_1 U10226 ( .ip(addr_resp[27]), .op(n9495) );
  mux2_1 U10227 ( .ip1(n9495), .ip2(addr_resp[27]), .s(n9494), .op(n9496) );
  nand4_1 U10228 ( .ip1(n9499), .ip2(n9498), .ip3(n9497), .ip4(n9496), .op(
        n9539) );
  inv_1 U10229 ( .ip(addr_resp[16]), .op(n9501) );
  mux2_1 U10230 ( .ip1(n9501), .ip2(addr_resp[16]), .s(n9500), .op(n9511) );
  inv_1 U10231 ( .ip(addr_resp[23]), .op(n9503) );
  mux2_1 U10232 ( .ip1(n9503), .ip2(addr_resp[23]), .s(n9502), .op(n9510) );
  inv_1 U10233 ( .ip(addr_resp[31]), .op(n9505) );
  mux2_1 U10234 ( .ip1(n9505), .ip2(addr_resp[31]), .s(n9504), .op(n9509) );
  inv_1 U10235 ( .ip(addr_resp[11]), .op(n9507) );
  mux2_1 U10236 ( .ip1(n9507), .ip2(addr_resp[11]), .s(n9506), .op(n9508) );
  nand4_1 U10237 ( .ip1(n9511), .ip2(n9510), .ip3(n9509), .ip4(n9508), .op(
        n9538) );
  inv_1 U10238 ( .ip(addr_resp[10]), .op(n9513) );
  mux2_1 U10239 ( .ip1(n9513), .ip2(addr_resp[10]), .s(n9512), .op(n9523) );
  inv_1 U10240 ( .ip(addr_resp[29]), .op(n9515) );
  mux2_1 U10241 ( .ip1(n9515), .ip2(addr_resp[29]), .s(n9514), .op(n9522) );
  inv_1 U10242 ( .ip(addr_resp[20]), .op(n9517) );
  mux2_1 U10243 ( .ip1(n9517), .ip2(addr_resp[20]), .s(n9516), .op(n9521) );
  inv_1 U10244 ( .ip(addr_resp[22]), .op(n9519) );
  mux2_1 U10245 ( .ip1(n9519), .ip2(addr_resp[22]), .s(n9518), .op(n9520) );
  nand4_1 U10246 ( .ip1(n9523), .ip2(n9522), .ip3(n9521), .ip4(n9520), .op(
        n9537) );
  inv_1 U10247 ( .ip(addr_resp[17]), .op(n9525) );
  mux2_1 U10248 ( .ip1(n9525), .ip2(addr_resp[17]), .s(n9524), .op(n9535) );
  inv_1 U10249 ( .ip(addr_resp[9]), .op(n9527) );
  mux2_1 U10250 ( .ip1(n9527), .ip2(addr_resp[9]), .s(n9526), .op(n9534) );
  inv_1 U10251 ( .ip(addr_resp[13]), .op(n9529) );
  mux2_1 U10252 ( .ip1(n9529), .ip2(addr_resp[13]), .s(n9528), .op(n9533) );
  inv_1 U10253 ( .ip(addr_resp[7]), .op(n9531) );
  mux2_1 U10254 ( .ip1(n9531), .ip2(addr_resp[7]), .s(n9530), .op(n9532) );
  nand4_1 U10255 ( .ip1(n9535), .ip2(n9534), .ip3(n9533), .ip4(n9532), .op(
        n9536) );
  nor4_1 U10256 ( .ip1(n9539), .ip2(n9538), .ip3(n9537), .ip4(n9536), .op(
        n9540) );
  nand4_1 U10257 ( .ip1(n9543), .ip2(n9542), .ip3(n9541), .ip4(n9540), .op(
        n9885) );
  inv_1 U10258 ( .ip(n9885), .op(n9925) );
  nor2_1 U10259 ( .ip1(n9544), .ip2(rd_temp), .op(n9846) );
  and2_1 U10260 ( .ip1(n9925), .ip2(n9846), .op(n9859) );
  nand2_1 U10261 ( .ip1(n9687), .ip2(n9859), .op(n9545) );
  nand2_1 U10262 ( .ip1(n9546), .ip2(n9545), .op(n9675) );
  nand2_1 U10263 ( .ip1(n9708), .ip2(n9675), .op(n9589) );
  mux2_1 U10264 ( .ip1(n9838), .ip2(\cache_data_A[0][25] ), .s(n9589), .op(
        n7384) );
  nand2_1 U10265 ( .ip1(data_rd_mem[26]), .ip2(n13295), .op(n9548) );
  nand2_1 U10266 ( .ip1(iCache_data_wr[26]), .ip2(n13294), .op(n9547) );
  nand2_1 U10267 ( .ip1(n9548), .ip2(n9547), .op(n9839) );
  mux2_1 U10268 ( .ip1(n9839), .ip2(\cache_data_A[0][26] ), .s(n9589), .op(
        n7383) );
  nand2_1 U10269 ( .ip1(data_rd_mem[27]), .ip2(n13295), .op(n9550) );
  nand2_1 U10270 ( .ip1(iCache_data_wr[27]), .ip2(n13294), .op(n9549) );
  nand2_1 U10271 ( .ip1(n9550), .ip2(n9549), .op(n9840) );
  mux2_1 U10272 ( .ip1(n9840), .ip2(\cache_data_A[0][27] ), .s(n9589), .op(
        n7382) );
  nand2_1 U10273 ( .ip1(data_rd_mem[28]), .ip2(n13295), .op(n9552) );
  nand2_1 U10274 ( .ip1(iCache_data_wr[28]), .ip2(n13294), .op(n9551) );
  nand2_1 U10275 ( .ip1(n9552), .ip2(n9551), .op(n9841) );
  mux2_1 U10276 ( .ip1(n9841), .ip2(\cache_data_A[0][28] ), .s(n9589), .op(
        n7381) );
  nand2_1 U10277 ( .ip1(data_rd_mem[29]), .ip2(n13295), .op(n9554) );
  nand2_1 U10278 ( .ip1(iCache_data_wr[29]), .ip2(n13294), .op(n9553) );
  nand2_1 U10279 ( .ip1(n9554), .ip2(n9553), .op(n9842) );
  mux2_1 U10280 ( .ip1(n9842), .ip2(\cache_data_A[0][29] ), .s(n9589), .op(
        n7380) );
  nand2_1 U10281 ( .ip1(data_rd_mem[30]), .ip2(n13295), .op(n9556) );
  nand2_1 U10282 ( .ip1(iCache_data_wr[30]), .ip2(n13294), .op(n9555) );
  nand2_1 U10283 ( .ip1(n9556), .ip2(n9555), .op(n9843) );
  mux2_1 U10284 ( .ip1(n9843), .ip2(\cache_data_A[0][30] ), .s(n9589), .op(
        n7379) );
  nand2_1 U10285 ( .ip1(data_rd_mem[31]), .ip2(n13295), .op(n9558) );
  nand2_1 U10286 ( .ip1(iCache_data_wr[31]), .ip2(n13294), .op(n9557) );
  nand2_1 U10287 ( .ip1(n9558), .ip2(n9557), .op(n9845) );
  mux2_1 U10288 ( .ip1(n9845), .ip2(\cache_data_A[0][31] ), .s(n9589), .op(
        n7378) );
  nand2_1 U10289 ( .ip1(data_rd_mem[0]), .ip2(n13295), .op(n9560) );
  nand2_1 U10290 ( .ip1(iCache_data_wr[0]), .ip2(n13294), .op(n9559) );
  nand2_1 U10291 ( .ip1(n9560), .ip2(n9559), .op(n9812) );
  mux2_1 U10292 ( .ip1(n9812), .ip2(\cache_data_A[0][0] ), .s(n9589), .op(
        n7377) );
  nand2_1 U10293 ( .ip1(data_rd_mem[1]), .ip2(n13295), .op(n9562) );
  nand2_1 U10294 ( .ip1(iCache_data_wr[1]), .ip2(n13294), .op(n9561) );
  nand2_1 U10295 ( .ip1(n9562), .ip2(n9561), .op(n9813) );
  mux2_1 U10296 ( .ip1(n9813), .ip2(\cache_data_A[0][1] ), .s(n9589), .op(
        n7376) );
  nand2_1 U10297 ( .ip1(data_rd_mem[2]), .ip2(n13295), .op(n9564) );
  nand2_1 U10298 ( .ip1(iCache_data_wr[2]), .ip2(n13294), .op(n9563) );
  nand2_1 U10299 ( .ip1(n9564), .ip2(n9563), .op(n9814) );
  mux2_1 U10300 ( .ip1(n9814), .ip2(\cache_data_A[0][2] ), .s(n9589), .op(
        n7375) );
  nand2_1 U10301 ( .ip1(data_rd_mem[3]), .ip2(n13295), .op(n9566) );
  nand2_1 U10302 ( .ip1(iCache_data_wr[3]), .ip2(n13294), .op(n9565) );
  nand2_1 U10303 ( .ip1(n9566), .ip2(n9565), .op(n9815) );
  buf_1 U10304 ( .ip(n9589), .op(n9610) );
  mux2_1 U10305 ( .ip1(n9815), .ip2(\cache_data_A[0][3] ), .s(n9610), .op(
        n7374) );
  nand2_1 U10306 ( .ip1(data_rd_mem[4]), .ip2(n13295), .op(n9568) );
  nand2_1 U10307 ( .ip1(iCache_data_wr[4]), .ip2(n9872), .op(n9567) );
  nand2_1 U10308 ( .ip1(n9568), .ip2(n9567), .op(n9816) );
  mux2_1 U10309 ( .ip1(n9816), .ip2(\cache_data_A[0][4] ), .s(n9589), .op(
        n7373) );
  nand2_1 U10310 ( .ip1(data_rd_mem[5]), .ip2(n13295), .op(n9570) );
  nand2_1 U10311 ( .ip1(iCache_data_wr[5]), .ip2(n13294), .op(n9569) );
  nand2_1 U10312 ( .ip1(n9570), .ip2(n9569), .op(n9817) );
  mux2_1 U10313 ( .ip1(n9817), .ip2(\cache_data_A[0][5] ), .s(n9589), .op(
        n7372) );
  nand2_1 U10314 ( .ip1(data_rd_mem[6]), .ip2(n13295), .op(n9572) );
  nand2_1 U10315 ( .ip1(iCache_data_wr[6]), .ip2(n13294), .op(n9571) );
  nand2_1 U10316 ( .ip1(n9572), .ip2(n9571), .op(n9818) );
  mux2_1 U10317 ( .ip1(n9818), .ip2(\cache_data_A[0][6] ), .s(n9589), .op(
        n7371) );
  nand2_1 U10318 ( .ip1(data_rd_mem[7]), .ip2(n13295), .op(n9574) );
  nand2_1 U10319 ( .ip1(iCache_data_wr[7]), .ip2(n13294), .op(n9573) );
  nand2_1 U10320 ( .ip1(n9574), .ip2(n9573), .op(n9819) );
  mux2_1 U10321 ( .ip1(n9819), .ip2(\cache_data_A[0][7] ), .s(n9589), .op(
        n7370) );
  nand2_1 U10322 ( .ip1(data_rd_mem[8]), .ip2(n13295), .op(n9576) );
  nand2_1 U10323 ( .ip1(iCache_data_wr[8]), .ip2(n13294), .op(n9575) );
  nand2_1 U10324 ( .ip1(n9576), .ip2(n9575), .op(n9820) );
  mux2_1 U10325 ( .ip1(n9820), .ip2(\cache_data_A[0][8] ), .s(n9589), .op(
        n7369) );
  nand2_1 U10326 ( .ip1(data_rd_mem[9]), .ip2(n13295), .op(n9578) );
  nand2_1 U10327 ( .ip1(iCache_data_wr[9]), .ip2(n13294), .op(n9577) );
  nand2_1 U10328 ( .ip1(n9578), .ip2(n9577), .op(n9821) );
  mux2_1 U10329 ( .ip1(n9821), .ip2(\cache_data_A[0][9] ), .s(n9589), .op(
        n7368) );
  nand2_1 U10330 ( .ip1(data_rd_mem[10]), .ip2(n13295), .op(n9580) );
  nand2_1 U10331 ( .ip1(iCache_data_wr[10]), .ip2(n13294), .op(n9579) );
  nand2_1 U10332 ( .ip1(n9580), .ip2(n9579), .op(n9822) );
  mux2_1 U10333 ( .ip1(n9822), .ip2(\cache_data_A[0][10] ), .s(n9589), .op(
        n7367) );
  nand2_1 U10334 ( .ip1(data_rd_mem[11]), .ip2(n13295), .op(n9582) );
  nand2_1 U10335 ( .ip1(iCache_data_wr[11]), .ip2(n13294), .op(n9581) );
  nand2_1 U10336 ( .ip1(n9582), .ip2(n9581), .op(n9823) );
  mux2_1 U10337 ( .ip1(n9823), .ip2(\cache_data_A[0][11] ), .s(n9589), .op(
        n7366) );
  nand2_1 U10338 ( .ip1(data_rd_mem[12]), .ip2(n13295), .op(n9584) );
  nand2_1 U10339 ( .ip1(iCache_data_wr[12]), .ip2(n13294), .op(n9583) );
  nand2_1 U10340 ( .ip1(n9584), .ip2(n9583), .op(n9824) );
  mux2_1 U10341 ( .ip1(n9824), .ip2(\cache_data_A[0][12] ), .s(n9589), .op(
        n7365) );
  nand2_1 U10342 ( .ip1(data_rd_mem[13]), .ip2(n13295), .op(n9586) );
  nand2_1 U10343 ( .ip1(iCache_data_wr[13]), .ip2(n13294), .op(n9585) );
  nand2_1 U10344 ( .ip1(n9586), .ip2(n9585), .op(n9825) );
  mux2_1 U10345 ( .ip1(n9825), .ip2(\cache_data_A[0][13] ), .s(n9589), .op(
        n7364) );
  nand2_1 U10346 ( .ip1(data_rd_mem[14]), .ip2(n13295), .op(n9588) );
  nand2_1 U10347 ( .ip1(iCache_data_wr[14]), .ip2(n13294), .op(n9587) );
  nand2_1 U10348 ( .ip1(n9588), .ip2(n9587), .op(n9826) );
  mux2_1 U10349 ( .ip1(n9826), .ip2(\cache_data_A[0][14] ), .s(n9589), .op(
        n7363) );
  nand2_1 U10350 ( .ip1(data_rd_mem[15]), .ip2(n13295), .op(n9591) );
  nand2_1 U10351 ( .ip1(iCache_data_wr[15]), .ip2(n13294), .op(n9590) );
  nand2_1 U10352 ( .ip1(n9591), .ip2(n9590), .op(n9827) );
  mux2_1 U10353 ( .ip1(n9827), .ip2(\cache_data_A[0][15] ), .s(n9610), .op(
        n7362) );
  nand2_1 U10354 ( .ip1(data_rd_mem[16]), .ip2(n13295), .op(n9593) );
  nand2_1 U10355 ( .ip1(iCache_data_wr[16]), .ip2(n13294), .op(n9592) );
  nand2_1 U10356 ( .ip1(n9593), .ip2(n9592), .op(n9828) );
  mux2_1 U10357 ( .ip1(n9828), .ip2(\cache_data_A[0][16] ), .s(n9610), .op(
        n7361) );
  nand2_1 U10358 ( .ip1(data_rd_mem[17]), .ip2(n13295), .op(n9595) );
  nand2_1 U10359 ( .ip1(iCache_data_wr[17]), .ip2(n13294), .op(n9594) );
  nand2_1 U10360 ( .ip1(n9595), .ip2(n9594), .op(n9829) );
  mux2_1 U10361 ( .ip1(n9829), .ip2(\cache_data_A[0][17] ), .s(n9610), .op(
        n7360) );
  nand2_1 U10362 ( .ip1(data_rd_mem[18]), .ip2(n13295), .op(n9597) );
  nand2_1 U10363 ( .ip1(iCache_data_wr[18]), .ip2(n9872), .op(n9596) );
  nand2_1 U10364 ( .ip1(n9597), .ip2(n9596), .op(n9830) );
  mux2_1 U10365 ( .ip1(n9830), .ip2(\cache_data_A[0][18] ), .s(n9610), .op(
        n7359) );
  nand2_1 U10366 ( .ip1(data_rd_mem[19]), .ip2(n13295), .op(n9599) );
  nand2_1 U10367 ( .ip1(iCache_data_wr[19]), .ip2(n9872), .op(n9598) );
  nand2_1 U10368 ( .ip1(n9599), .ip2(n9598), .op(n9831) );
  mux2_1 U10369 ( .ip1(n9831), .ip2(\cache_data_A[0][19] ), .s(n9610), .op(
        n7358) );
  nand2_1 U10370 ( .ip1(data_rd_mem[20]), .ip2(n13295), .op(n9601) );
  nand2_1 U10371 ( .ip1(iCache_data_wr[20]), .ip2(n9872), .op(n9600) );
  nand2_1 U10372 ( .ip1(n9601), .ip2(n9600), .op(n9832) );
  mux2_1 U10373 ( .ip1(n9832), .ip2(\cache_data_A[0][20] ), .s(n9610), .op(
        n7357) );
  nand2_1 U10374 ( .ip1(data_rd_mem[21]), .ip2(n13295), .op(n9603) );
  nand2_1 U10375 ( .ip1(iCache_data_wr[21]), .ip2(n9872), .op(n9602) );
  nand2_1 U10376 ( .ip1(n9603), .ip2(n9602), .op(n9833) );
  mux2_1 U10377 ( .ip1(n9833), .ip2(\cache_data_A[0][21] ), .s(n9610), .op(
        n7356) );
  nand2_1 U10378 ( .ip1(data_rd_mem[22]), .ip2(n13295), .op(n9605) );
  nand2_1 U10379 ( .ip1(iCache_data_wr[22]), .ip2(n9872), .op(n9604) );
  nand2_1 U10380 ( .ip1(n9605), .ip2(n9604), .op(n9835) );
  mux2_1 U10381 ( .ip1(n9835), .ip2(\cache_data_A[0][22] ), .s(n9610), .op(
        n7355) );
  nand2_1 U10382 ( .ip1(data_rd_mem[23]), .ip2(n13295), .op(n9607) );
  nand2_1 U10383 ( .ip1(iCache_data_wr[23]), .ip2(n9872), .op(n9606) );
  nand2_1 U10384 ( .ip1(n9607), .ip2(n9606), .op(n9836) );
  mux2_1 U10385 ( .ip1(n9836), .ip2(\cache_data_A[0][23] ), .s(n9610), .op(
        n7354) );
  nand2_1 U10386 ( .ip1(data_rd_mem[24]), .ip2(n13295), .op(n9609) );
  nand2_1 U10387 ( .ip1(iCache_data_wr[24]), .ip2(n9872), .op(n9608) );
  nand2_1 U10388 ( .ip1(n9609), .ip2(n9608), .op(n9837) );
  mux2_1 U10389 ( .ip1(n9837), .ip2(\cache_data_A[0][24] ), .s(n9610), .op(
        n7353) );
  nor3_1 U10390 ( .ip1(SelectWay), .ip2(mem_data_cnt[3]), .ip3(n9700), .op(
        n13162) );
  nand2_1 U10391 ( .ip1(n13162), .ip2(n9619), .op(n9612) );
  nor3_1 U10392 ( .ip1(addr_resp[3]), .ip2(n9705), .ip3(n9885), .op(n12595) );
  nand2_1 U10393 ( .ip1(n12595), .ip2(n9846), .op(n9611) );
  nand2_1 U10394 ( .ip1(n9612), .ip2(n9611), .op(n9678) );
  nand2_1 U10395 ( .ip1(n9708), .ip2(n9678), .op(n9613) );
  mux2_1 U10396 ( .ip1(n9812), .ip2(\cache_data_A[0][32] ), .s(n9613), .op(
        n7352) );
  mux2_1 U10397 ( .ip1(n9813), .ip2(\cache_data_A[0][33] ), .s(n9613), .op(
        n7351) );
  mux2_1 U10398 ( .ip1(n9814), .ip2(\cache_data_A[0][34] ), .s(n9613), .op(
        n7350) );
  mux2_1 U10399 ( .ip1(n9815), .ip2(\cache_data_A[0][35] ), .s(n9613), .op(
        n7349) );
  mux2_1 U10400 ( .ip1(n9816), .ip2(\cache_data_A[0][36] ), .s(n9613), .op(
        n7348) );
  mux2_1 U10401 ( .ip1(n9817), .ip2(\cache_data_A[0][37] ), .s(n9613), .op(
        n7347) );
  mux2_1 U10402 ( .ip1(n9818), .ip2(\cache_data_A[0][38] ), .s(n9613), .op(
        n7346) );
  mux2_1 U10403 ( .ip1(n9819), .ip2(\cache_data_A[0][39] ), .s(n9613), .op(
        n7345) );
  mux2_1 U10404 ( .ip1(n9820), .ip2(\cache_data_A[0][40] ), .s(n9613), .op(
        n7344) );
  mux2_1 U10405 ( .ip1(n9821), .ip2(\cache_data_A[0][41] ), .s(n9613), .op(
        n7343) );
  buf_1 U10406 ( .ip(n9613), .op(n9614) );
  mux2_1 U10407 ( .ip1(n9822), .ip2(\cache_data_A[0][42] ), .s(n9614), .op(
        n7342) );
  mux2_1 U10408 ( .ip1(n9823), .ip2(\cache_data_A[0][43] ), .s(n9613), .op(
        n7341) );
  mux2_1 U10409 ( .ip1(n9824), .ip2(\cache_data_A[0][44] ), .s(n9613), .op(
        n7340) );
  mux2_1 U10410 ( .ip1(n9825), .ip2(\cache_data_A[0][45] ), .s(n9613), .op(
        n7339) );
  mux2_1 U10411 ( .ip1(n9826), .ip2(\cache_data_A[0][46] ), .s(n9613), .op(
        n7338) );
  mux2_1 U10412 ( .ip1(n9827), .ip2(\cache_data_A[0][47] ), .s(n9613), .op(
        n7337) );
  mux2_1 U10413 ( .ip1(n9828), .ip2(\cache_data_A[0][48] ), .s(n9614), .op(
        n7336) );
  mux2_1 U10414 ( .ip1(n9829), .ip2(\cache_data_A[0][49] ), .s(n9614), .op(
        n7335) );
  mux2_1 U10415 ( .ip1(n9830), .ip2(\cache_data_A[0][50] ), .s(n9614), .op(
        n7334) );
  mux2_1 U10416 ( .ip1(n9831), .ip2(\cache_data_A[0][51] ), .s(n9613), .op(
        n7333) );
  mux2_1 U10417 ( .ip1(n9832), .ip2(\cache_data_A[0][52] ), .s(n9613), .op(
        n7332) );
  mux2_1 U10418 ( .ip1(n9833), .ip2(\cache_data_A[0][53] ), .s(n9613), .op(
        n7331) );
  mux2_1 U10419 ( .ip1(n9835), .ip2(\cache_data_A[0][54] ), .s(n9613), .op(
        n7330) );
  mux2_1 U10420 ( .ip1(n9836), .ip2(\cache_data_A[0][55] ), .s(n9613), .op(
        n7329) );
  mux2_1 U10421 ( .ip1(n9837), .ip2(\cache_data_A[0][56] ), .s(n9613), .op(
        n7328) );
  mux2_1 U10422 ( .ip1(n9838), .ip2(\cache_data_A[0][57] ), .s(n9614), .op(
        n7327) );
  mux2_1 U10423 ( .ip1(n9839), .ip2(\cache_data_A[0][58] ), .s(n9614), .op(
        n7326) );
  mux2_1 U10424 ( .ip1(n9840), .ip2(\cache_data_A[0][59] ), .s(n9614), .op(
        n7325) );
  mux2_1 U10425 ( .ip1(n9841), .ip2(\cache_data_A[0][60] ), .s(n9614), .op(
        n7324) );
  mux2_1 U10426 ( .ip1(n9842), .ip2(\cache_data_A[0][61] ), .s(n9614), .op(
        n7323) );
  mux2_1 U10427 ( .ip1(n9843), .ip2(\cache_data_A[0][62] ), .s(n9614), .op(
        n7322) );
  mux2_1 U10428 ( .ip1(n9845), .ip2(\cache_data_A[0][63] ), .s(n9614), .op(
        n7321) );
  buf_1 U10429 ( .ip(n9812), .op(n9770) );
  nand3_1 U10430 ( .ip1(n9702), .ip2(n9700), .ip3(mem_data_cnt[3]), .op(n13163) );
  or2_1 U10431 ( .ip1(n13163), .ip2(n13191), .op(n9616) );
  nor2_1 U10432 ( .ip1(addr_resp[2]), .ip2(n9704), .op(n9905) );
  nand2_1 U10433 ( .ip1(n9859), .ip2(n9905), .op(n9615) );
  nand2_1 U10434 ( .ip1(n9616), .ip2(n9615), .op(n9660) );
  nand2_1 U10435 ( .ip1(n13293), .ip2(n9660), .op(n9681) );
  nor2_1 U10436 ( .ip1(n9860), .ip2(n9681), .op(n9617) );
  mux2_1 U10437 ( .ip1(\cache_data_A[0][64] ), .ip2(n9770), .s(n9617), .op(
        n7320) );
  mux2_1 U10438 ( .ip1(\cache_data_A[0][65] ), .ip2(n9813), .s(n9617), .op(
        n7319) );
  mux2_1 U10439 ( .ip1(\cache_data_A[0][66] ), .ip2(n9814), .s(n9617), .op(
        n7318) );
  mux2_1 U10440 ( .ip1(\cache_data_A[0][67] ), .ip2(n9815), .s(n9617), .op(
        n7317) );
  mux2_1 U10441 ( .ip1(\cache_data_A[0][68] ), .ip2(n9816), .s(n9617), .op(
        n7316) );
  mux2_1 U10442 ( .ip1(\cache_data_A[0][69] ), .ip2(n9817), .s(n9617), .op(
        n7315) );
  mux2_1 U10443 ( .ip1(\cache_data_A[0][70] ), .ip2(n9818), .s(n9617), .op(
        n7314) );
  mux2_1 U10444 ( .ip1(\cache_data_A[0][71] ), .ip2(n9819), .s(n9617), .op(
        n7313) );
  mux2_1 U10445 ( .ip1(\cache_data_A[0][72] ), .ip2(n9820), .s(n9617), .op(
        n7312) );
  buf_1 U10446 ( .ip(n9617), .op(n9618) );
  mux2_1 U10447 ( .ip1(\cache_data_A[0][73] ), .ip2(n9821), .s(n9618), .op(
        n7311) );
  mux2_1 U10448 ( .ip1(\cache_data_A[0][74] ), .ip2(n9822), .s(n9618), .op(
        n7310) );
  mux2_1 U10449 ( .ip1(\cache_data_A[0][75] ), .ip2(n9823), .s(n9617), .op(
        n7309) );
  mux2_1 U10450 ( .ip1(\cache_data_A[0][76] ), .ip2(n9824), .s(n9617), .op(
        n7308) );
  mux2_1 U10451 ( .ip1(\cache_data_A[0][77] ), .ip2(n9825), .s(n9618), .op(
        n7307) );
  mux2_1 U10452 ( .ip1(\cache_data_A[0][78] ), .ip2(n9826), .s(n9617), .op(
        n7306) );
  mux2_1 U10453 ( .ip1(\cache_data_A[0][79] ), .ip2(n9827), .s(n9617), .op(
        n7305) );
  mux2_1 U10454 ( .ip1(\cache_data_A[0][80] ), .ip2(n9828), .s(n9617), .op(
        n7304) );
  buf_1 U10455 ( .ip(n9829), .op(n9787) );
  mux2_1 U10456 ( .ip1(\cache_data_A[0][81] ), .ip2(n9787), .s(n9617), .op(
        n7303) );
  buf_1 U10457 ( .ip(n9830), .op(n9788) );
  mux2_1 U10458 ( .ip1(\cache_data_A[0][82] ), .ip2(n9788), .s(n9617), .op(
        n7302) );
  mux2_1 U10459 ( .ip1(\cache_data_A[0][83] ), .ip2(n9831), .s(n9617), .op(
        n7301) );
  mux2_1 U10460 ( .ip1(\cache_data_A[0][84] ), .ip2(n9832), .s(n9617), .op(
        n7300) );
  mux2_1 U10461 ( .ip1(\cache_data_A[0][85] ), .ip2(n9833), .s(n9617), .op(
        n7299) );
  mux2_1 U10462 ( .ip1(\cache_data_A[0][86] ), .ip2(n9835), .s(n9617), .op(
        n7298) );
  mux2_1 U10463 ( .ip1(\cache_data_A[0][87] ), .ip2(n9836), .s(n9617), .op(
        n7297) );
  mux2_1 U10464 ( .ip1(\cache_data_A[0][88] ), .ip2(n9837), .s(n9618), .op(
        n7296) );
  buf_1 U10465 ( .ip(n9838), .op(n9796) );
  mux2_1 U10466 ( .ip1(\cache_data_A[0][89] ), .ip2(n9796), .s(n9618), .op(
        n7295) );
  buf_1 U10467 ( .ip(n9839), .op(n9797) );
  mux2_1 U10468 ( .ip1(\cache_data_A[0][90] ), .ip2(n9797), .s(n9618), .op(
        n7294) );
  buf_1 U10469 ( .ip(n9840), .op(n9798) );
  mux2_1 U10470 ( .ip1(\cache_data_A[0][91] ), .ip2(n9798), .s(n9618), .op(
        n7293) );
  buf_1 U10471 ( .ip(n9841), .op(n9799) );
  mux2_1 U10472 ( .ip1(\cache_data_A[0][92] ), .ip2(n9799), .s(n9618), .op(
        n7292) );
  buf_1 U10473 ( .ip(n9842), .op(n9800) );
  mux2_1 U10474 ( .ip1(\cache_data_A[0][93] ), .ip2(n9800), .s(n9618), .op(
        n7291) );
  buf_1 U10475 ( .ip(n9843), .op(n9801) );
  mux2_1 U10476 ( .ip1(\cache_data_A[0][94] ), .ip2(n9801), .s(n9618), .op(
        n7290) );
  buf_1 U10477 ( .ip(n9845), .op(n9803) );
  mux2_1 U10478 ( .ip1(\cache_data_A[0][95] ), .ip2(n9803), .s(n9618), .op(
        n7289) );
  nor3_1 U10479 ( .ip1(SelectWay), .ip2(n9701), .ip3(n9700), .op(n13172) );
  nand2_1 U10480 ( .ip1(n13172), .ip2(n9619), .op(n9621) );
  nor3_1 U10481 ( .ip1(n9704), .ip2(n9705), .ip3(n9885), .op(n12509) );
  nand2_1 U10482 ( .ip1(n12509), .ip2(n9846), .op(n9620) );
  nand2_1 U10483 ( .ip1(n9621), .ip2(n9620), .op(n9684) );
  nand2_1 U10484 ( .ip1(n9708), .ip2(n9684), .op(n9622) );
  mux2_1 U10485 ( .ip1(n9799), .ip2(\cache_data_A[0][124] ), .s(n9622), .op(
        n7288) );
  mux2_1 U10486 ( .ip1(n9800), .ip2(\cache_data_A[0][125] ), .s(n9622), .op(
        n7287) );
  mux2_1 U10487 ( .ip1(n9801), .ip2(\cache_data_A[0][126] ), .s(n9622), .op(
        n7286) );
  mux2_1 U10488 ( .ip1(n9803), .ip2(\cache_data_A[0][127] ), .s(n9622), .op(
        n7285) );
  mux2_1 U10489 ( .ip1(n9770), .ip2(\cache_data_A[0][96] ), .s(n9622), .op(
        n7284) );
  buf_1 U10490 ( .ip(n9813), .op(n9771) );
  mux2_1 U10491 ( .ip1(n9771), .ip2(\cache_data_A[0][97] ), .s(n9622), .op(
        n7283) );
  buf_1 U10492 ( .ip(n9814), .op(n9772) );
  mux2_1 U10493 ( .ip1(n9772), .ip2(\cache_data_A[0][98] ), .s(n9622), .op(
        n7282) );
  buf_1 U10494 ( .ip(n9815), .op(n9773) );
  mux2_1 U10495 ( .ip1(n9773), .ip2(\cache_data_A[0][99] ), .s(n9622), .op(
        n7281) );
  buf_1 U10496 ( .ip(n9816), .op(n9774) );
  mux2_1 U10497 ( .ip1(n9774), .ip2(\cache_data_A[0][100] ), .s(n9622), .op(
        n7280) );
  buf_1 U10498 ( .ip(n9817), .op(n9775) );
  mux2_1 U10499 ( .ip1(n9775), .ip2(\cache_data_A[0][101] ), .s(n9622), .op(
        n7279) );
  buf_1 U10500 ( .ip(n9818), .op(n9776) );
  mux2_1 U10501 ( .ip1(n9776), .ip2(\cache_data_A[0][102] ), .s(n9622), .op(
        n7278) );
  buf_1 U10502 ( .ip(n9819), .op(n9777) );
  mux2_1 U10503 ( .ip1(n9777), .ip2(\cache_data_A[0][103] ), .s(n9622), .op(
        n7277) );
  buf_1 U10504 ( .ip(n9820), .op(n9778) );
  mux2_1 U10505 ( .ip1(n9778), .ip2(\cache_data_A[0][104] ), .s(n9622), .op(
        n7276) );
  buf_1 U10506 ( .ip(n9821), .op(n9779) );
  mux2_1 U10507 ( .ip1(n9779), .ip2(\cache_data_A[0][105] ), .s(n9622), .op(
        n7275) );
  buf_1 U10508 ( .ip(n9822), .op(n9780) );
  mux2_1 U10509 ( .ip1(n9780), .ip2(\cache_data_A[0][106] ), .s(n9622), .op(
        n7274) );
  buf_1 U10510 ( .ip(n9823), .op(n9781) );
  mux2_1 U10511 ( .ip1(n9781), .ip2(\cache_data_A[0][107] ), .s(n9622), .op(
        n7273) );
  buf_1 U10512 ( .ip(n9824), .op(n9782) );
  mux2_1 U10513 ( .ip1(n9782), .ip2(\cache_data_A[0][108] ), .s(n9622), .op(
        n7272) );
  buf_1 U10514 ( .ip(n9825), .op(n9783) );
  mux2_1 U10515 ( .ip1(n9783), .ip2(\cache_data_A[0][109] ), .s(n9622), .op(
        n7271) );
  buf_1 U10516 ( .ip(n9826), .op(n9784) );
  buf_1 U10517 ( .ip(n9622), .op(n9623) );
  mux2_1 U10518 ( .ip1(n9784), .ip2(\cache_data_A[0][110] ), .s(n9623), .op(
        n7270) );
  buf_1 U10519 ( .ip(n9827), .op(n9785) );
  mux2_1 U10520 ( .ip1(n9785), .ip2(\cache_data_A[0][111] ), .s(n9623), .op(
        n7269) );
  buf_1 U10521 ( .ip(n9828), .op(n9786) );
  mux2_1 U10522 ( .ip1(n9786), .ip2(\cache_data_A[0][112] ), .s(n9622), .op(
        n7268) );
  mux2_1 U10523 ( .ip1(n9787), .ip2(\cache_data_A[0][113] ), .s(n9623), .op(
        n7267) );
  mux2_1 U10524 ( .ip1(n9788), .ip2(\cache_data_A[0][114] ), .s(n9623), .op(
        n7266) );
  buf_1 U10525 ( .ip(n9831), .op(n9789) );
  mux2_1 U10526 ( .ip1(n9789), .ip2(\cache_data_A[0][115] ), .s(n9623), .op(
        n7265) );
  buf_1 U10527 ( .ip(n9832), .op(n9790) );
  mux2_1 U10528 ( .ip1(n9790), .ip2(\cache_data_A[0][116] ), .s(n9622), .op(
        n7264) );
  buf_1 U10529 ( .ip(n9833), .op(n9791) );
  mux2_1 U10530 ( .ip1(n9791), .ip2(\cache_data_A[0][117] ), .s(n9622), .op(
        n7263) );
  buf_1 U10531 ( .ip(n9835), .op(n9792) );
  mux2_1 U10532 ( .ip1(n9792), .ip2(\cache_data_A[0][118] ), .s(n9623), .op(
        n7262) );
  buf_1 U10533 ( .ip(n9836), .op(n9794) );
  mux2_1 U10534 ( .ip1(n9794), .ip2(\cache_data_A[0][119] ), .s(n9623), .op(
        n7261) );
  buf_1 U10535 ( .ip(n9837), .op(n9795) );
  mux2_1 U10536 ( .ip1(n9795), .ip2(\cache_data_A[0][120] ), .s(n9623), .op(
        n7260) );
  mux2_1 U10537 ( .ip1(n9796), .ip2(\cache_data_A[0][121] ), .s(n9623), .op(
        n7259) );
  mux2_1 U10538 ( .ip1(n9797), .ip2(\cache_data_A[0][122] ), .s(n9623), .op(
        n7258) );
  mux2_1 U10539 ( .ip1(n9798), .ip2(\cache_data_A[0][123] ), .s(n9623), .op(
        n7257) );
  nand2_1 U10540 ( .ip1(n13293), .ip2(n9675), .op(n9665) );
  nor2_1 U10541 ( .ip1(n9862), .ip2(n9665), .op(n9624) );
  mux2_1 U10542 ( .ip1(\cache_data_A[1][0] ), .ip2(n9812), .s(n9624), .op(
        n7256) );
  mux2_1 U10543 ( .ip1(\cache_data_A[1][1] ), .ip2(n9813), .s(n9624), .op(
        n7255) );
  mux2_1 U10544 ( .ip1(\cache_data_A[1][2] ), .ip2(n9814), .s(n9624), .op(
        n7254) );
  mux2_1 U10545 ( .ip1(\cache_data_A[1][3] ), .ip2(n9815), .s(n9624), .op(
        n7253) );
  mux2_1 U10546 ( .ip1(\cache_data_A[1][4] ), .ip2(n9816), .s(n9624), .op(
        n7252) );
  mux2_1 U10547 ( .ip1(\cache_data_A[1][5] ), .ip2(n9817), .s(n9624), .op(
        n7251) );
  mux2_1 U10548 ( .ip1(\cache_data_A[1][6] ), .ip2(n9818), .s(n9624), .op(
        n7250) );
  mux2_1 U10549 ( .ip1(\cache_data_A[1][7] ), .ip2(n9819), .s(n9624), .op(
        n7249) );
  mux2_1 U10550 ( .ip1(\cache_data_A[1][8] ), .ip2(n9820), .s(n9624), .op(
        n7248) );
  buf_1 U10551 ( .ip(n9624), .op(n9625) );
  mux2_1 U10552 ( .ip1(\cache_data_A[1][9] ), .ip2(n9821), .s(n9625), .op(
        n7247) );
  mux2_1 U10553 ( .ip1(\cache_data_A[1][10] ), .ip2(n9822), .s(n9625), .op(
        n7246) );
  mux2_1 U10554 ( .ip1(\cache_data_A[1][11] ), .ip2(n9823), .s(n9624), .op(
        n7245) );
  mux2_1 U10555 ( .ip1(\cache_data_A[1][12] ), .ip2(n9824), .s(n9624), .op(
        n7244) );
  mux2_1 U10556 ( .ip1(\cache_data_A[1][13] ), .ip2(n9825), .s(n9625), .op(
        n7243) );
  mux2_1 U10557 ( .ip1(\cache_data_A[1][14] ), .ip2(n9826), .s(n9624), .op(
        n7242) );
  mux2_1 U10558 ( .ip1(\cache_data_A[1][15] ), .ip2(n9827), .s(n9624), .op(
        n7241) );
  mux2_1 U10559 ( .ip1(\cache_data_A[1][16] ), .ip2(n9828), .s(n9624), .op(
        n7240) );
  mux2_1 U10560 ( .ip1(\cache_data_A[1][17] ), .ip2(n9829), .s(n9624), .op(
        n7239) );
  mux2_1 U10561 ( .ip1(\cache_data_A[1][18] ), .ip2(n9830), .s(n9624), .op(
        n7238) );
  mux2_1 U10562 ( .ip1(\cache_data_A[1][19] ), .ip2(n9831), .s(n9624), .op(
        n7237) );
  mux2_1 U10563 ( .ip1(\cache_data_A[1][20] ), .ip2(n9832), .s(n9624), .op(
        n7236) );
  mux2_1 U10564 ( .ip1(\cache_data_A[1][21] ), .ip2(n9833), .s(n9624), .op(
        n7235) );
  mux2_1 U10565 ( .ip1(\cache_data_A[1][22] ), .ip2(n9835), .s(n9624), .op(
        n7234) );
  mux2_1 U10566 ( .ip1(\cache_data_A[1][23] ), .ip2(n9836), .s(n9624), .op(
        n7233) );
  mux2_1 U10567 ( .ip1(\cache_data_A[1][24] ), .ip2(n9837), .s(n9625), .op(
        n7232) );
  mux2_1 U10568 ( .ip1(\cache_data_A[1][25] ), .ip2(n9838), .s(n9625), .op(
        n7231) );
  mux2_1 U10569 ( .ip1(\cache_data_A[1][26] ), .ip2(n9839), .s(n9625), .op(
        n7230) );
  mux2_1 U10570 ( .ip1(\cache_data_A[1][27] ), .ip2(n9840), .s(n9625), .op(
        n7229) );
  mux2_1 U10571 ( .ip1(\cache_data_A[1][28] ), .ip2(n9841), .s(n9625), .op(
        n7228) );
  mux2_1 U10572 ( .ip1(\cache_data_A[1][29] ), .ip2(n9842), .s(n9625), .op(
        n7227) );
  mux2_1 U10573 ( .ip1(\cache_data_A[1][30] ), .ip2(n9843), .s(n9625), .op(
        n7226) );
  mux2_1 U10574 ( .ip1(\cache_data_A[1][31] ), .ip2(n9845), .s(n9625), .op(
        n7225) );
  nand2_1 U10575 ( .ip1(n9717), .ip2(n9678), .op(n9626) );
  mux2_1 U10576 ( .ip1(n9812), .ip2(\cache_data_A[1][32] ), .s(n9626), .op(
        n7224) );
  mux2_1 U10577 ( .ip1(n9813), .ip2(\cache_data_A[1][33] ), .s(n9626), .op(
        n7223) );
  mux2_1 U10578 ( .ip1(n9814), .ip2(\cache_data_A[1][34] ), .s(n9626), .op(
        n7222) );
  mux2_1 U10579 ( .ip1(n9815), .ip2(\cache_data_A[1][35] ), .s(n9626), .op(
        n7221) );
  mux2_1 U10580 ( .ip1(n9816), .ip2(\cache_data_A[1][36] ), .s(n9626), .op(
        n7220) );
  mux2_1 U10581 ( .ip1(n9817), .ip2(\cache_data_A[1][37] ), .s(n9626), .op(
        n7219) );
  mux2_1 U10582 ( .ip1(n9818), .ip2(\cache_data_A[1][38] ), .s(n9626), .op(
        n7218) );
  mux2_1 U10583 ( .ip1(n9819), .ip2(\cache_data_A[1][39] ), .s(n9626), .op(
        n7217) );
  mux2_1 U10584 ( .ip1(n9820), .ip2(\cache_data_A[1][40] ), .s(n9626), .op(
        n7216) );
  buf_1 U10585 ( .ip(n9626), .op(n9627) );
  mux2_1 U10586 ( .ip1(n9821), .ip2(\cache_data_A[1][41] ), .s(n9627), .op(
        n7215) );
  mux2_1 U10587 ( .ip1(n9822), .ip2(\cache_data_A[1][42] ), .s(n9626), .op(
        n7214) );
  mux2_1 U10588 ( .ip1(n9823), .ip2(\cache_data_A[1][43] ), .s(n9626), .op(
        n7213) );
  mux2_1 U10589 ( .ip1(n9824), .ip2(\cache_data_A[1][44] ), .s(n9626), .op(
        n7212) );
  mux2_1 U10590 ( .ip1(n9825), .ip2(\cache_data_A[1][45] ), .s(n9626), .op(
        n7211) );
  mux2_1 U10591 ( .ip1(n9826), .ip2(\cache_data_A[1][46] ), .s(n9626), .op(
        n7210) );
  mux2_1 U10592 ( .ip1(n9827), .ip2(\cache_data_A[1][47] ), .s(n9626), .op(
        n7209) );
  mux2_1 U10593 ( .ip1(n9828), .ip2(\cache_data_A[1][48] ), .s(n9626), .op(
        n7208) );
  mux2_1 U10594 ( .ip1(n9829), .ip2(\cache_data_A[1][49] ), .s(n9626), .op(
        n7207) );
  mux2_1 U10595 ( .ip1(n9830), .ip2(\cache_data_A[1][50] ), .s(n9626), .op(
        n7206) );
  mux2_1 U10596 ( .ip1(n9831), .ip2(\cache_data_A[1][51] ), .s(n9626), .op(
        n7205) );
  mux2_1 U10597 ( .ip1(n9790), .ip2(\cache_data_A[1][52] ), .s(n9626), .op(
        n7204) );
  mux2_1 U10598 ( .ip1(n9833), .ip2(\cache_data_A[1][53] ), .s(n9626), .op(
        n7203) );
  mux2_1 U10599 ( .ip1(n9835), .ip2(\cache_data_A[1][54] ), .s(n9627), .op(
        n7202) );
  mux2_1 U10600 ( .ip1(n9836), .ip2(\cache_data_A[1][55] ), .s(n9627), .op(
        n7201) );
  mux2_1 U10601 ( .ip1(n9837), .ip2(\cache_data_A[1][56] ), .s(n9627), .op(
        n7200) );
  mux2_1 U10602 ( .ip1(n9838), .ip2(\cache_data_A[1][57] ), .s(n9627), .op(
        n7199) );
  mux2_1 U10603 ( .ip1(n9839), .ip2(\cache_data_A[1][58] ), .s(n9627), .op(
        n7198) );
  mux2_1 U10604 ( .ip1(n9840), .ip2(\cache_data_A[1][59] ), .s(n9627), .op(
        n7197) );
  mux2_1 U10605 ( .ip1(n9841), .ip2(\cache_data_A[1][60] ), .s(n9627), .op(
        n7196) );
  mux2_1 U10606 ( .ip1(n9842), .ip2(\cache_data_A[1][61] ), .s(n9627), .op(
        n7195) );
  mux2_1 U10607 ( .ip1(n9843), .ip2(\cache_data_A[1][62] ), .s(n9627), .op(
        n7194) );
  mux2_1 U10608 ( .ip1(n9845), .ip2(\cache_data_A[1][63] ), .s(n9627), .op(
        n7193) );
  nand2_1 U10609 ( .ip1(n9717), .ip2(n9660), .op(n9628) );
  mux2_1 U10610 ( .ip1(n9845), .ip2(\cache_data_A[1][95] ), .s(n9628), .op(
        n7192) );
  mux2_1 U10611 ( .ip1(n9812), .ip2(\cache_data_A[1][64] ), .s(n9628), .op(
        n7191) );
  mux2_1 U10612 ( .ip1(n9813), .ip2(\cache_data_A[1][65] ), .s(n9628), .op(
        n7190) );
  mux2_1 U10613 ( .ip1(n9814), .ip2(\cache_data_A[1][66] ), .s(n9628), .op(
        n7189) );
  mux2_1 U10614 ( .ip1(n9815), .ip2(\cache_data_A[1][67] ), .s(n9628), .op(
        n7188) );
  mux2_1 U10615 ( .ip1(n9816), .ip2(\cache_data_A[1][68] ), .s(n9628), .op(
        n7187) );
  mux2_1 U10616 ( .ip1(n9817), .ip2(\cache_data_A[1][69] ), .s(n9628), .op(
        n7186) );
  mux2_1 U10617 ( .ip1(n9818), .ip2(\cache_data_A[1][70] ), .s(n9628), .op(
        n7185) );
  mux2_1 U10618 ( .ip1(n9819), .ip2(\cache_data_A[1][71] ), .s(n9628), .op(
        n7184) );
  buf_1 U10619 ( .ip(n9628), .op(n9629) );
  mux2_1 U10620 ( .ip1(n9820), .ip2(\cache_data_A[1][72] ), .s(n9629), .op(
        n7183) );
  mux2_1 U10621 ( .ip1(n9821), .ip2(\cache_data_A[1][73] ), .s(n9628), .op(
        n7182) );
  mux2_1 U10622 ( .ip1(n9822), .ip2(\cache_data_A[1][74] ), .s(n9628), .op(
        n7181) );
  mux2_1 U10623 ( .ip1(n9823), .ip2(\cache_data_A[1][75] ), .s(n9628), .op(
        n7180) );
  mux2_1 U10624 ( .ip1(n9824), .ip2(\cache_data_A[1][76] ), .s(n9628), .op(
        n7179) );
  mux2_1 U10625 ( .ip1(n9825), .ip2(\cache_data_A[1][77] ), .s(n9628), .op(
        n7178) );
  mux2_1 U10626 ( .ip1(n9826), .ip2(\cache_data_A[1][78] ), .s(n9628), .op(
        n7177) );
  mux2_1 U10627 ( .ip1(n9827), .ip2(\cache_data_A[1][79] ), .s(n9628), .op(
        n7176) );
  mux2_1 U10628 ( .ip1(n9828), .ip2(\cache_data_A[1][80] ), .s(n9628), .op(
        n7175) );
  mux2_1 U10629 ( .ip1(n9829), .ip2(\cache_data_A[1][81] ), .s(n9628), .op(
        n7174) );
  mux2_1 U10630 ( .ip1(n9830), .ip2(\cache_data_A[1][82] ), .s(n9628), .op(
        n7173) );
  mux2_1 U10631 ( .ip1(n9831), .ip2(\cache_data_A[1][83] ), .s(n9628), .op(
        n7172) );
  mux2_1 U10632 ( .ip1(n9832), .ip2(\cache_data_A[1][84] ), .s(n9628), .op(
        n7171) );
  mux2_1 U10633 ( .ip1(n9833), .ip2(\cache_data_A[1][85] ), .s(n9629), .op(
        n7170) );
  mux2_1 U10634 ( .ip1(n9835), .ip2(\cache_data_A[1][86] ), .s(n9629), .op(
        n7169) );
  mux2_1 U10635 ( .ip1(n9836), .ip2(\cache_data_A[1][87] ), .s(n9629), .op(
        n7168) );
  mux2_1 U10636 ( .ip1(n9837), .ip2(\cache_data_A[1][88] ), .s(n9629), .op(
        n7167) );
  mux2_1 U10637 ( .ip1(n9838), .ip2(\cache_data_A[1][89] ), .s(n9629), .op(
        n7166) );
  mux2_1 U10638 ( .ip1(n9839), .ip2(\cache_data_A[1][90] ), .s(n9629), .op(
        n7165) );
  mux2_1 U10639 ( .ip1(n9840), .ip2(\cache_data_A[1][91] ), .s(n9629), .op(
        n7164) );
  mux2_1 U10640 ( .ip1(n9841), .ip2(\cache_data_A[1][92] ), .s(n9629), .op(
        n7163) );
  mux2_1 U10641 ( .ip1(n9842), .ip2(\cache_data_A[1][93] ), .s(n9629), .op(
        n7162) );
  mux2_1 U10642 ( .ip1(n9843), .ip2(\cache_data_A[1][94] ), .s(n9629), .op(
        n7161) );
  nand2_1 U10643 ( .ip1(n13293), .ip2(n9684), .op(n9672) );
  nor2_1 U10644 ( .ip1(n9862), .ip2(n9672), .op(n9630) );
  mux2_1 U10645 ( .ip1(\cache_data_A[1][96] ), .ip2(n9770), .s(n9630), .op(
        n7160) );
  mux2_1 U10646 ( .ip1(\cache_data_A[1][97] ), .ip2(n9813), .s(n9630), .op(
        n7159) );
  mux2_1 U10647 ( .ip1(\cache_data_A[1][98] ), .ip2(n9814), .s(n9630), .op(
        n7158) );
  mux2_1 U10648 ( .ip1(\cache_data_A[1][99] ), .ip2(n9815), .s(n9630), .op(
        n7157) );
  mux2_1 U10649 ( .ip1(\cache_data_A[1][100] ), .ip2(n9816), .s(n9630), .op(
        n7156) );
  mux2_1 U10650 ( .ip1(\cache_data_A[1][101] ), .ip2(n9817), .s(n9630), .op(
        n7155) );
  mux2_1 U10651 ( .ip1(\cache_data_A[1][102] ), .ip2(n9818), .s(n9630), .op(
        n7154) );
  mux2_1 U10652 ( .ip1(\cache_data_A[1][103] ), .ip2(n9819), .s(n9630), .op(
        n7153) );
  mux2_1 U10653 ( .ip1(\cache_data_A[1][104] ), .ip2(n9820), .s(n9630), .op(
        n7152) );
  buf_1 U10654 ( .ip(n9630), .op(n9631) );
  mux2_1 U10655 ( .ip1(\cache_data_A[1][105] ), .ip2(n9821), .s(n9631), .op(
        n7151) );
  mux2_1 U10656 ( .ip1(\cache_data_A[1][106] ), .ip2(n9822), .s(n9631), .op(
        n7150) );
  mux2_1 U10657 ( .ip1(\cache_data_A[1][107] ), .ip2(n9823), .s(n9630), .op(
        n7149) );
  mux2_1 U10658 ( .ip1(\cache_data_A[1][108] ), .ip2(n9824), .s(n9630), .op(
        n7148) );
  mux2_1 U10659 ( .ip1(\cache_data_A[1][109] ), .ip2(n9825), .s(n9631), .op(
        n7147) );
  mux2_1 U10660 ( .ip1(\cache_data_A[1][110] ), .ip2(n9826), .s(n9630), .op(
        n7146) );
  mux2_1 U10661 ( .ip1(\cache_data_A[1][111] ), .ip2(n9827), .s(n9630), .op(
        n7145) );
  mux2_1 U10662 ( .ip1(\cache_data_A[1][112] ), .ip2(n9828), .s(n9630), .op(
        n7144) );
  mux2_1 U10663 ( .ip1(\cache_data_A[1][113] ), .ip2(n9787), .s(n9630), .op(
        n7143) );
  mux2_1 U10664 ( .ip1(\cache_data_A[1][114] ), .ip2(n9788), .s(n9630), .op(
        n7142) );
  mux2_1 U10665 ( .ip1(\cache_data_A[1][115] ), .ip2(n9831), .s(n9630), .op(
        n7141) );
  mux2_1 U10666 ( .ip1(\cache_data_A[1][116] ), .ip2(n9832), .s(n9630), .op(
        n7140) );
  mux2_1 U10667 ( .ip1(\cache_data_A[1][117] ), .ip2(n9833), .s(n9630), .op(
        n7139) );
  mux2_1 U10668 ( .ip1(\cache_data_A[1][118] ), .ip2(n9835), .s(n9630), .op(
        n7138) );
  mux2_1 U10669 ( .ip1(\cache_data_A[1][119] ), .ip2(n9836), .s(n9630), .op(
        n7137) );
  mux2_1 U10670 ( .ip1(\cache_data_A[1][120] ), .ip2(n9837), .s(n9631), .op(
        n7136) );
  mux2_1 U10671 ( .ip1(\cache_data_A[1][121] ), .ip2(n9796), .s(n9631), .op(
        n7135) );
  mux2_1 U10672 ( .ip1(\cache_data_A[1][122] ), .ip2(n9797), .s(n9631), .op(
        n7134) );
  mux2_1 U10673 ( .ip1(\cache_data_A[1][123] ), .ip2(n9798), .s(n9631), .op(
        n7133) );
  mux2_1 U10674 ( .ip1(\cache_data_A[1][124] ), .ip2(n9799), .s(n9631), .op(
        n7132) );
  mux2_1 U10675 ( .ip1(\cache_data_A[1][125] ), .ip2(n9800), .s(n9631), .op(
        n7131) );
  mux2_1 U10676 ( .ip1(\cache_data_A[1][126] ), .ip2(n9801), .s(n9631), .op(
        n7130) );
  mux2_1 U10677 ( .ip1(\cache_data_A[1][127] ), .ip2(n9803), .s(n9631), .op(
        n7129) );
  nor2_1 U10678 ( .ip1(n9864), .ip2(n9665), .op(n9632) );
  mux2_1 U10679 ( .ip1(\cache_data_A[2][0] ), .ip2(n9812), .s(n9632), .op(
        n7128) );
  mux2_1 U10680 ( .ip1(\cache_data_A[2][1] ), .ip2(n9771), .s(n9632), .op(
        n7127) );
  mux2_1 U10681 ( .ip1(\cache_data_A[2][2] ), .ip2(n9772), .s(n9632), .op(
        n7126) );
  mux2_1 U10682 ( .ip1(\cache_data_A[2][3] ), .ip2(n9773), .s(n9632), .op(
        n7125) );
  mux2_1 U10683 ( .ip1(\cache_data_A[2][4] ), .ip2(n9774), .s(n9632), .op(
        n7124) );
  mux2_1 U10684 ( .ip1(\cache_data_A[2][5] ), .ip2(n9775), .s(n9632), .op(
        n7123) );
  mux2_1 U10685 ( .ip1(\cache_data_A[2][6] ), .ip2(n9776), .s(n9632), .op(
        n7122) );
  mux2_1 U10686 ( .ip1(\cache_data_A[2][7] ), .ip2(n9777), .s(n9632), .op(
        n7121) );
  mux2_1 U10687 ( .ip1(\cache_data_A[2][8] ), .ip2(n9778), .s(n9632), .op(
        n7120) );
  buf_1 U10688 ( .ip(n9632), .op(n9633) );
  mux2_1 U10689 ( .ip1(\cache_data_A[2][9] ), .ip2(n9779), .s(n9633), .op(
        n7119) );
  mux2_1 U10690 ( .ip1(\cache_data_A[2][10] ), .ip2(n9780), .s(n9633), .op(
        n7118) );
  mux2_1 U10691 ( .ip1(\cache_data_A[2][11] ), .ip2(n9781), .s(n9632), .op(
        n7117) );
  mux2_1 U10692 ( .ip1(\cache_data_A[2][12] ), .ip2(n9782), .s(n9632), .op(
        n7116) );
  mux2_1 U10693 ( .ip1(\cache_data_A[2][13] ), .ip2(n9783), .s(n9633), .op(
        n7115) );
  mux2_1 U10694 ( .ip1(\cache_data_A[2][14] ), .ip2(n9784), .s(n9632), .op(
        n7114) );
  mux2_1 U10695 ( .ip1(\cache_data_A[2][15] ), .ip2(n9785), .s(n9632), .op(
        n7113) );
  mux2_1 U10696 ( .ip1(\cache_data_A[2][16] ), .ip2(n9786), .s(n9632), .op(
        n7112) );
  mux2_1 U10697 ( .ip1(\cache_data_A[2][17] ), .ip2(n9829), .s(n9632), .op(
        n7111) );
  mux2_1 U10698 ( .ip1(\cache_data_A[2][18] ), .ip2(n9830), .s(n9632), .op(
        n7110) );
  mux2_1 U10699 ( .ip1(\cache_data_A[2][19] ), .ip2(n9831), .s(n9632), .op(
        n7109) );
  mux2_1 U10700 ( .ip1(\cache_data_A[2][20] ), .ip2(n9832), .s(n9632), .op(
        n7108) );
  mux2_1 U10701 ( .ip1(\cache_data_A[2][21] ), .ip2(n9833), .s(n9632), .op(
        n7107) );
  mux2_1 U10702 ( .ip1(\cache_data_A[2][22] ), .ip2(n9835), .s(n9632), .op(
        n7106) );
  mux2_1 U10703 ( .ip1(\cache_data_A[2][23] ), .ip2(n9836), .s(n9632), .op(
        n7105) );
  mux2_1 U10704 ( .ip1(\cache_data_A[2][24] ), .ip2(n9837), .s(n9633), .op(
        n7104) );
  mux2_1 U10705 ( .ip1(\cache_data_A[2][25] ), .ip2(n9838), .s(n9633), .op(
        n7103) );
  mux2_1 U10706 ( .ip1(\cache_data_A[2][26] ), .ip2(n9839), .s(n9633), .op(
        n7102) );
  mux2_1 U10707 ( .ip1(\cache_data_A[2][27] ), .ip2(n9840), .s(n9633), .op(
        n7101) );
  mux2_1 U10708 ( .ip1(\cache_data_A[2][28] ), .ip2(n9841), .s(n9633), .op(
        n7100) );
  mux2_1 U10709 ( .ip1(\cache_data_A[2][29] ), .ip2(n9842), .s(n9633), .op(
        n7099) );
  mux2_1 U10710 ( .ip1(\cache_data_A[2][30] ), .ip2(n9843), .s(n9633), .op(
        n7098) );
  mux2_1 U10711 ( .ip1(\cache_data_A[2][31] ), .ip2(n9845), .s(n9633), .op(
        n7097) );
  nand2_1 U10712 ( .ip1(n9726), .ip2(n9678), .op(n9634) );
  mux2_1 U10713 ( .ip1(n9812), .ip2(\cache_data_A[2][32] ), .s(n9634), .op(
        n7096) );
  mux2_1 U10714 ( .ip1(n9813), .ip2(\cache_data_A[2][33] ), .s(n9634), .op(
        n7095) );
  mux2_1 U10715 ( .ip1(n9814), .ip2(\cache_data_A[2][34] ), .s(n9634), .op(
        n7094) );
  mux2_1 U10716 ( .ip1(n9815), .ip2(\cache_data_A[2][35] ), .s(n9634), .op(
        n7093) );
  mux2_1 U10717 ( .ip1(n9816), .ip2(\cache_data_A[2][36] ), .s(n9634), .op(
        n7092) );
  mux2_1 U10718 ( .ip1(n9817), .ip2(\cache_data_A[2][37] ), .s(n9634), .op(
        n7091) );
  mux2_1 U10719 ( .ip1(n9818), .ip2(\cache_data_A[2][38] ), .s(n9634), .op(
        n7090) );
  mux2_1 U10720 ( .ip1(n9819), .ip2(\cache_data_A[2][39] ), .s(n9634), .op(
        n7089) );
  mux2_1 U10721 ( .ip1(n9820), .ip2(\cache_data_A[2][40] ), .s(n9634), .op(
        n7088) );
  mux2_1 U10722 ( .ip1(n9821), .ip2(\cache_data_A[2][41] ), .s(n9634), .op(
        n7087) );
  mux2_1 U10723 ( .ip1(n9822), .ip2(\cache_data_A[2][42] ), .s(n9634), .op(
        n7086) );
  mux2_1 U10724 ( .ip1(n9823), .ip2(\cache_data_A[2][43] ), .s(n9634), .op(
        n7085) );
  buf_1 U10725 ( .ip(n9634), .op(n9635) );
  mux2_1 U10726 ( .ip1(n9824), .ip2(\cache_data_A[2][44] ), .s(n9635), .op(
        n7084) );
  mux2_1 U10727 ( .ip1(n9825), .ip2(\cache_data_A[2][45] ), .s(n9634), .op(
        n7083) );
  mux2_1 U10728 ( .ip1(n9826), .ip2(\cache_data_A[2][46] ), .s(n9634), .op(
        n7082) );
  mux2_1 U10729 ( .ip1(n9827), .ip2(\cache_data_A[2][47] ), .s(n9634), .op(
        n7081) );
  mux2_1 U10730 ( .ip1(n9828), .ip2(\cache_data_A[2][48] ), .s(n9635), .op(
        n7080) );
  mux2_1 U10731 ( .ip1(n9829), .ip2(\cache_data_A[2][49] ), .s(n9634), .op(
        n7079) );
  mux2_1 U10732 ( .ip1(n9830), .ip2(\cache_data_A[2][50] ), .s(n9634), .op(
        n7078) );
  mux2_1 U10733 ( .ip1(n9831), .ip2(\cache_data_A[2][51] ), .s(n9634), .op(
        n7077) );
  mux2_1 U10734 ( .ip1(n9832), .ip2(\cache_data_A[2][52] ), .s(n9634), .op(
        n7076) );
  mux2_1 U10735 ( .ip1(n9833), .ip2(\cache_data_A[2][53] ), .s(n9634), .op(
        n7075) );
  mux2_1 U10736 ( .ip1(n9835), .ip2(\cache_data_A[2][54] ), .s(n9634), .op(
        n7074) );
  mux2_1 U10737 ( .ip1(n9836), .ip2(\cache_data_A[2][55] ), .s(n9635), .op(
        n7073) );
  mux2_1 U10738 ( .ip1(n9837), .ip2(\cache_data_A[2][56] ), .s(n9635), .op(
        n7072) );
  mux2_1 U10739 ( .ip1(n9838), .ip2(\cache_data_A[2][57] ), .s(n9635), .op(
        n7071) );
  mux2_1 U10740 ( .ip1(n9839), .ip2(\cache_data_A[2][58] ), .s(n9635), .op(
        n7070) );
  mux2_1 U10741 ( .ip1(n9840), .ip2(\cache_data_A[2][59] ), .s(n9635), .op(
        n7069) );
  mux2_1 U10742 ( .ip1(n9841), .ip2(\cache_data_A[2][60] ), .s(n9635), .op(
        n7068) );
  mux2_1 U10743 ( .ip1(n9842), .ip2(\cache_data_A[2][61] ), .s(n9635), .op(
        n7067) );
  mux2_1 U10744 ( .ip1(n9843), .ip2(\cache_data_A[2][62] ), .s(n9635), .op(
        n7066) );
  mux2_1 U10745 ( .ip1(n9845), .ip2(\cache_data_A[2][63] ), .s(n9635), .op(
        n7065) );
  nand2_1 U10746 ( .ip1(n9726), .ip2(n9660), .op(n9636) );
  mux2_1 U10747 ( .ip1(n9772), .ip2(\cache_data_A[2][66] ), .s(n9636), .op(
        n7064) );
  mux2_1 U10748 ( .ip1(n9773), .ip2(\cache_data_A[2][67] ), .s(n9636), .op(
        n7063) );
  mux2_1 U10749 ( .ip1(n9774), .ip2(\cache_data_A[2][68] ), .s(n9636), .op(
        n7062) );
  mux2_1 U10750 ( .ip1(n9775), .ip2(\cache_data_A[2][69] ), .s(n9636), .op(
        n7061) );
  mux2_1 U10751 ( .ip1(n9776), .ip2(\cache_data_A[2][70] ), .s(n9636), .op(
        n7060) );
  mux2_1 U10752 ( .ip1(n9777), .ip2(\cache_data_A[2][71] ), .s(n9636), .op(
        n7059) );
  mux2_1 U10753 ( .ip1(n9778), .ip2(\cache_data_A[2][72] ), .s(n9636), .op(
        n7058) );
  mux2_1 U10754 ( .ip1(n9779), .ip2(\cache_data_A[2][73] ), .s(n9636), .op(
        n7057) );
  mux2_1 U10755 ( .ip1(n9780), .ip2(\cache_data_A[2][74] ), .s(n9636), .op(
        n7056) );
  buf_1 U10756 ( .ip(n9636), .op(n9637) );
  mux2_1 U10757 ( .ip1(n9781), .ip2(\cache_data_A[2][75] ), .s(n9637), .op(
        n7055) );
  mux2_1 U10758 ( .ip1(n9782), .ip2(\cache_data_A[2][76] ), .s(n9636), .op(
        n7054) );
  mux2_1 U10759 ( .ip1(n9783), .ip2(\cache_data_A[2][77] ), .s(n9636), .op(
        n7053) );
  mux2_1 U10760 ( .ip1(n9784), .ip2(\cache_data_A[2][78] ), .s(n9636), .op(
        n7052) );
  mux2_1 U10761 ( .ip1(n9785), .ip2(\cache_data_A[2][79] ), .s(n9636), .op(
        n7051) );
  mux2_1 U10762 ( .ip1(n9786), .ip2(\cache_data_A[2][80] ), .s(n9636), .op(
        n7050) );
  mux2_1 U10763 ( .ip1(n9787), .ip2(\cache_data_A[2][81] ), .s(n9636), .op(
        n7049) );
  mux2_1 U10764 ( .ip1(n9788), .ip2(\cache_data_A[2][82] ), .s(n9636), .op(
        n7048) );
  mux2_1 U10765 ( .ip1(n9789), .ip2(\cache_data_A[2][83] ), .s(n9636), .op(
        n7047) );
  mux2_1 U10766 ( .ip1(n9790), .ip2(\cache_data_A[2][84] ), .s(n9636), .op(
        n7046) );
  mux2_1 U10767 ( .ip1(n9791), .ip2(\cache_data_A[2][85] ), .s(n9636), .op(
        n7045) );
  mux2_1 U10768 ( .ip1(n9792), .ip2(\cache_data_A[2][86] ), .s(n9636), .op(
        n7044) );
  mux2_1 U10769 ( .ip1(n9794), .ip2(\cache_data_A[2][87] ), .s(n9636), .op(
        n7043) );
  mux2_1 U10770 ( .ip1(n9795), .ip2(\cache_data_A[2][88] ), .s(n9637), .op(
        n7042) );
  mux2_1 U10771 ( .ip1(n9796), .ip2(\cache_data_A[2][89] ), .s(n9637), .op(
        n7041) );
  mux2_1 U10772 ( .ip1(n9797), .ip2(\cache_data_A[2][90] ), .s(n9637), .op(
        n7040) );
  mux2_1 U10773 ( .ip1(n9798), .ip2(\cache_data_A[2][91] ), .s(n9637), .op(
        n7039) );
  mux2_1 U10774 ( .ip1(n9799), .ip2(\cache_data_A[2][92] ), .s(n9637), .op(
        n7038) );
  mux2_1 U10775 ( .ip1(n9800), .ip2(\cache_data_A[2][93] ), .s(n9637), .op(
        n7037) );
  mux2_1 U10776 ( .ip1(n9801), .ip2(\cache_data_A[2][94] ), .s(n9637), .op(
        n7036) );
  mux2_1 U10777 ( .ip1(n9803), .ip2(\cache_data_A[2][95] ), .s(n9637), .op(
        n7035) );
  mux2_1 U10778 ( .ip1(n9770), .ip2(\cache_data_A[2][64] ), .s(n9637), .op(
        n7034) );
  mux2_1 U10779 ( .ip1(n9771), .ip2(\cache_data_A[2][65] ), .s(n9637), .op(
        n7033) );
  nor2_1 U10780 ( .ip1(n9864), .ip2(n9672), .op(n9638) );
  mux2_1 U10781 ( .ip1(\cache_data_A[2][96] ), .ip2(n9770), .s(n9638), .op(
        n7032) );
  mux2_1 U10782 ( .ip1(\cache_data_A[2][97] ), .ip2(n9771), .s(n9638), .op(
        n7031) );
  mux2_1 U10783 ( .ip1(\cache_data_A[2][98] ), .ip2(n9772), .s(n9638), .op(
        n7030) );
  mux2_1 U10784 ( .ip1(\cache_data_A[2][99] ), .ip2(n9773), .s(n9638), .op(
        n7029) );
  mux2_1 U10785 ( .ip1(\cache_data_A[2][100] ), .ip2(n9774), .s(n9638), .op(
        n7028) );
  mux2_1 U10786 ( .ip1(\cache_data_A[2][101] ), .ip2(n9775), .s(n9638), .op(
        n7027) );
  mux2_1 U10787 ( .ip1(\cache_data_A[2][102] ), .ip2(n9776), .s(n9638), .op(
        n7026) );
  mux2_1 U10788 ( .ip1(\cache_data_A[2][103] ), .ip2(n9777), .s(n9638), .op(
        n7025) );
  mux2_1 U10789 ( .ip1(\cache_data_A[2][104] ), .ip2(n9778), .s(n9638), .op(
        n7024) );
  buf_1 U10790 ( .ip(n9638), .op(n9639) );
  mux2_1 U10791 ( .ip1(\cache_data_A[2][105] ), .ip2(n9779), .s(n9639), .op(
        n7023) );
  mux2_1 U10792 ( .ip1(\cache_data_A[2][106] ), .ip2(n9780), .s(n9639), .op(
        n7022) );
  mux2_1 U10793 ( .ip1(\cache_data_A[2][107] ), .ip2(n9781), .s(n9638), .op(
        n7021) );
  mux2_1 U10794 ( .ip1(\cache_data_A[2][108] ), .ip2(n9782), .s(n9638), .op(
        n7020) );
  mux2_1 U10795 ( .ip1(\cache_data_A[2][109] ), .ip2(n9783), .s(n9639), .op(
        n7019) );
  mux2_1 U10796 ( .ip1(\cache_data_A[2][110] ), .ip2(n9784), .s(n9638), .op(
        n7018) );
  mux2_1 U10797 ( .ip1(\cache_data_A[2][111] ), .ip2(n9785), .s(n9638), .op(
        n7017) );
  mux2_1 U10798 ( .ip1(\cache_data_A[2][112] ), .ip2(n9786), .s(n9638), .op(
        n7016) );
  mux2_1 U10799 ( .ip1(\cache_data_A[2][113] ), .ip2(n9787), .s(n9638), .op(
        n7015) );
  mux2_1 U10800 ( .ip1(\cache_data_A[2][114] ), .ip2(n9788), .s(n9638), .op(
        n7014) );
  mux2_1 U10801 ( .ip1(\cache_data_A[2][115] ), .ip2(n9831), .s(n9638), .op(
        n7013) );
  mux2_1 U10802 ( .ip1(\cache_data_A[2][116] ), .ip2(n9832), .s(n9638), .op(
        n7012) );
  mux2_1 U10803 ( .ip1(\cache_data_A[2][117] ), .ip2(n9833), .s(n9638), .op(
        n7011) );
  mux2_1 U10804 ( .ip1(\cache_data_A[2][118] ), .ip2(n9835), .s(n9638), .op(
        n7010) );
  mux2_1 U10805 ( .ip1(\cache_data_A[2][119] ), .ip2(n9836), .s(n9638), .op(
        n7009) );
  mux2_1 U10806 ( .ip1(\cache_data_A[2][120] ), .ip2(n9837), .s(n9639), .op(
        n7008) );
  mux2_1 U10807 ( .ip1(\cache_data_A[2][121] ), .ip2(n9796), .s(n9639), .op(
        n7007) );
  mux2_1 U10808 ( .ip1(\cache_data_A[2][122] ), .ip2(n9797), .s(n9639), .op(
        n7006) );
  mux2_1 U10809 ( .ip1(\cache_data_A[2][123] ), .ip2(n9798), .s(n9639), .op(
        n7005) );
  mux2_1 U10810 ( .ip1(\cache_data_A[2][124] ), .ip2(n9799), .s(n9639), .op(
        n7004) );
  mux2_1 U10811 ( .ip1(\cache_data_A[2][125] ), .ip2(n9800), .s(n9639), .op(
        n7003) );
  mux2_1 U10812 ( .ip1(\cache_data_A[2][126] ), .ip2(n9801), .s(n9639), .op(
        n7002) );
  mux2_1 U10813 ( .ip1(\cache_data_A[2][127] ), .ip2(n9803), .s(n9639), .op(
        n7001) );
  nor2_1 U10814 ( .ip1(n9866), .ip2(n9665), .op(n9640) );
  mux2_1 U10815 ( .ip1(\cache_data_A[3][0] ), .ip2(n9812), .s(n9640), .op(
        n7000) );
  mux2_1 U10816 ( .ip1(\cache_data_A[3][1] ), .ip2(n9813), .s(n9640), .op(
        n6999) );
  mux2_1 U10817 ( .ip1(\cache_data_A[3][2] ), .ip2(n9814), .s(n9640), .op(
        n6998) );
  mux2_1 U10818 ( .ip1(\cache_data_A[3][3] ), .ip2(n9815), .s(n9640), .op(
        n6997) );
  mux2_1 U10819 ( .ip1(\cache_data_A[3][4] ), .ip2(n9816), .s(n9640), .op(
        n6996) );
  mux2_1 U10820 ( .ip1(\cache_data_A[3][5] ), .ip2(n9817), .s(n9640), .op(
        n6995) );
  mux2_1 U10821 ( .ip1(\cache_data_A[3][6] ), .ip2(n9818), .s(n9640), .op(
        n6994) );
  mux2_1 U10822 ( .ip1(\cache_data_A[3][7] ), .ip2(n9819), .s(n9640), .op(
        n6993) );
  mux2_1 U10823 ( .ip1(\cache_data_A[3][8] ), .ip2(n9820), .s(n9640), .op(
        n6992) );
  mux2_1 U10824 ( .ip1(\cache_data_A[3][9] ), .ip2(n9821), .s(n9640), .op(
        n6991) );
  mux2_1 U10825 ( .ip1(\cache_data_A[3][10] ), .ip2(n9822), .s(n9640), .op(
        n6990) );
  mux2_1 U10826 ( .ip1(\cache_data_A[3][11] ), .ip2(n9823), .s(n9640), .op(
        n6989) );
  mux2_1 U10827 ( .ip1(\cache_data_A[3][12] ), .ip2(n9824), .s(n9640), .op(
        n6988) );
  mux2_1 U10828 ( .ip1(\cache_data_A[3][13] ), .ip2(n9825), .s(n9640), .op(
        n6987) );
  mux2_1 U10829 ( .ip1(\cache_data_A[3][14] ), .ip2(n9826), .s(n9640), .op(
        n6986) );
  mux2_1 U10830 ( .ip1(\cache_data_A[3][15] ), .ip2(n9827), .s(n9640), .op(
        n6985) );
  mux2_1 U10831 ( .ip1(\cache_data_A[3][16] ), .ip2(n9828), .s(n9640), .op(
        n6984) );
  mux2_1 U10832 ( .ip1(\cache_data_A[3][17] ), .ip2(n9829), .s(n9640), .op(
        n6983) );
  mux2_1 U10833 ( .ip1(\cache_data_A[3][18] ), .ip2(n9830), .s(n9640), .op(
        n6982) );
  buf_1 U10834 ( .ip(n9640), .op(n9641) );
  mux2_1 U10835 ( .ip1(\cache_data_A[3][19] ), .ip2(n9831), .s(n9641), .op(
        n6981) );
  mux2_1 U10836 ( .ip1(\cache_data_A[3][20] ), .ip2(n9832), .s(n9641), .op(
        n6980) );
  mux2_1 U10837 ( .ip1(\cache_data_A[3][21] ), .ip2(n9833), .s(n9641), .op(
        n6979) );
  mux2_1 U10838 ( .ip1(\cache_data_A[3][22] ), .ip2(n9835), .s(n9641), .op(
        n6978) );
  mux2_1 U10839 ( .ip1(\cache_data_A[3][23] ), .ip2(n9836), .s(n9641), .op(
        n6977) );
  mux2_1 U10840 ( .ip1(\cache_data_A[3][24] ), .ip2(n9837), .s(n9640), .op(
        n6976) );
  mux2_1 U10841 ( .ip1(\cache_data_A[3][25] ), .ip2(n9838), .s(n9640), .op(
        n6975) );
  mux2_1 U10842 ( .ip1(\cache_data_A[3][26] ), .ip2(n9839), .s(n9641), .op(
        n6974) );
  mux2_1 U10843 ( .ip1(\cache_data_A[3][27] ), .ip2(n9840), .s(n9641), .op(
        n6973) );
  mux2_1 U10844 ( .ip1(\cache_data_A[3][28] ), .ip2(n9841), .s(n9641), .op(
        n6972) );
  mux2_1 U10845 ( .ip1(\cache_data_A[3][29] ), .ip2(n9842), .s(n9641), .op(
        n6971) );
  mux2_1 U10846 ( .ip1(\cache_data_A[3][30] ), .ip2(n9843), .s(n9641), .op(
        n6970) );
  mux2_1 U10847 ( .ip1(\cache_data_A[3][31] ), .ip2(n9845), .s(n9641), .op(
        n6969) );
  nand2_1 U10848 ( .ip1(n9735), .ip2(n9678), .op(n9642) );
  mux2_1 U10849 ( .ip1(n9817), .ip2(\cache_data_A[3][37] ), .s(n9642), .op(
        n6968) );
  buf_1 U10850 ( .ip(n9642), .op(n9643) );
  mux2_1 U10851 ( .ip1(n9818), .ip2(\cache_data_A[3][38] ), .s(n9643), .op(
        n6967) );
  mux2_1 U10852 ( .ip1(n9819), .ip2(\cache_data_A[3][39] ), .s(n9642), .op(
        n6966) );
  mux2_1 U10853 ( .ip1(n9820), .ip2(\cache_data_A[3][40] ), .s(n9642), .op(
        n6965) );
  mux2_1 U10854 ( .ip1(n9821), .ip2(\cache_data_A[3][41] ), .s(n9642), .op(
        n6964) );
  mux2_1 U10855 ( .ip1(n9822), .ip2(\cache_data_A[3][42] ), .s(n9642), .op(
        n6963) );
  mux2_1 U10856 ( .ip1(n9823), .ip2(\cache_data_A[3][43] ), .s(n9642), .op(
        n6962) );
  mux2_1 U10857 ( .ip1(n9824), .ip2(\cache_data_A[3][44] ), .s(n9642), .op(
        n6961) );
  mux2_1 U10858 ( .ip1(n9825), .ip2(\cache_data_A[3][45] ), .s(n9642), .op(
        n6960) );
  mux2_1 U10859 ( .ip1(n9826), .ip2(\cache_data_A[3][46] ), .s(n9642), .op(
        n6959) );
  mux2_1 U10860 ( .ip1(n9827), .ip2(\cache_data_A[3][47] ), .s(n9642), .op(
        n6958) );
  mux2_1 U10861 ( .ip1(n9828), .ip2(\cache_data_A[3][48] ), .s(n9642), .op(
        n6957) );
  mux2_1 U10862 ( .ip1(n9829), .ip2(\cache_data_A[3][49] ), .s(n9642), .op(
        n6956) );
  mux2_1 U10863 ( .ip1(n9830), .ip2(\cache_data_A[3][50] ), .s(n9642), .op(
        n6955) );
  mux2_1 U10864 ( .ip1(n9831), .ip2(\cache_data_A[3][51] ), .s(n9643), .op(
        n6954) );
  mux2_1 U10865 ( .ip1(n9832), .ip2(\cache_data_A[3][52] ), .s(n9642), .op(
        n6953) );
  mux2_1 U10866 ( .ip1(n9833), .ip2(\cache_data_A[3][53] ), .s(n9642), .op(
        n6952) );
  mux2_1 U10867 ( .ip1(n9835), .ip2(\cache_data_A[3][54] ), .s(n9642), .op(
        n6951) );
  mux2_1 U10868 ( .ip1(n9836), .ip2(\cache_data_A[3][55] ), .s(n9642), .op(
        n6950) );
  mux2_1 U10869 ( .ip1(n9837), .ip2(\cache_data_A[3][56] ), .s(n9642), .op(
        n6949) );
  mux2_1 U10870 ( .ip1(n9838), .ip2(\cache_data_A[3][57] ), .s(n9642), .op(
        n6948) );
  mux2_1 U10871 ( .ip1(n9839), .ip2(\cache_data_A[3][58] ), .s(n9642), .op(
        n6947) );
  mux2_1 U10872 ( .ip1(n9840), .ip2(\cache_data_A[3][59] ), .s(n9642), .op(
        n6946) );
  mux2_1 U10873 ( .ip1(n9841), .ip2(\cache_data_A[3][60] ), .s(n9643), .op(
        n6945) );
  mux2_1 U10874 ( .ip1(n9842), .ip2(\cache_data_A[3][61] ), .s(n9643), .op(
        n6944) );
  mux2_1 U10875 ( .ip1(n9843), .ip2(\cache_data_A[3][62] ), .s(n9643), .op(
        n6943) );
  mux2_1 U10876 ( .ip1(n9845), .ip2(\cache_data_A[3][63] ), .s(n9643), .op(
        n6942) );
  mux2_1 U10877 ( .ip1(n9812), .ip2(\cache_data_A[3][32] ), .s(n9643), .op(
        n6941) );
  mux2_1 U10878 ( .ip1(n9813), .ip2(\cache_data_A[3][33] ), .s(n9643), .op(
        n6940) );
  mux2_1 U10879 ( .ip1(n9814), .ip2(\cache_data_A[3][34] ), .s(n9643), .op(
        n6939) );
  mux2_1 U10880 ( .ip1(n9815), .ip2(\cache_data_A[3][35] ), .s(n9643), .op(
        n6938) );
  mux2_1 U10881 ( .ip1(n9816), .ip2(\cache_data_A[3][36] ), .s(n9643), .op(
        n6937) );
  nor2_1 U10882 ( .ip1(n9866), .ip2(n9681), .op(n9644) );
  mux2_1 U10883 ( .ip1(\cache_data_A[3][64] ), .ip2(n9770), .s(n9644), .op(
        n6936) );
  mux2_1 U10884 ( .ip1(\cache_data_A[3][65] ), .ip2(n9771), .s(n9644), .op(
        n6935) );
  mux2_1 U10885 ( .ip1(\cache_data_A[3][66] ), .ip2(n9772), .s(n9644), .op(
        n6934) );
  mux2_1 U10886 ( .ip1(\cache_data_A[3][67] ), .ip2(n9773), .s(n9644), .op(
        n6933) );
  mux2_1 U10887 ( .ip1(\cache_data_A[3][68] ), .ip2(n9774), .s(n9644), .op(
        n6932) );
  mux2_1 U10888 ( .ip1(\cache_data_A[3][69] ), .ip2(n9775), .s(n9644), .op(
        n6931) );
  mux2_1 U10889 ( .ip1(\cache_data_A[3][70] ), .ip2(n9776), .s(n9644), .op(
        n6930) );
  mux2_1 U10890 ( .ip1(\cache_data_A[3][71] ), .ip2(n9777), .s(n9644), .op(
        n6929) );
  mux2_1 U10891 ( .ip1(\cache_data_A[3][72] ), .ip2(n9778), .s(n9644), .op(
        n6928) );
  mux2_1 U10892 ( .ip1(\cache_data_A[3][73] ), .ip2(n9779), .s(n9644), .op(
        n6927) );
  mux2_1 U10893 ( .ip1(\cache_data_A[3][74] ), .ip2(n9780), .s(n9644), .op(
        n6926) );
  mux2_1 U10894 ( .ip1(\cache_data_A[3][75] ), .ip2(n9781), .s(n9644), .op(
        n6925) );
  mux2_1 U10895 ( .ip1(\cache_data_A[3][76] ), .ip2(n9782), .s(n9644), .op(
        n6924) );
  mux2_1 U10896 ( .ip1(\cache_data_A[3][77] ), .ip2(n9783), .s(n9644), .op(
        n6923) );
  mux2_1 U10897 ( .ip1(\cache_data_A[3][78] ), .ip2(n9784), .s(n9644), .op(
        n6922) );
  mux2_1 U10898 ( .ip1(\cache_data_A[3][79] ), .ip2(n9785), .s(n9644), .op(
        n6921) );
  mux2_1 U10899 ( .ip1(\cache_data_A[3][80] ), .ip2(n9786), .s(n9644), .op(
        n6920) );
  mux2_1 U10900 ( .ip1(\cache_data_A[3][81] ), .ip2(n9787), .s(n9644), .op(
        n6919) );
  mux2_1 U10901 ( .ip1(\cache_data_A[3][82] ), .ip2(n9788), .s(n9644), .op(
        n6918) );
  buf_1 U10902 ( .ip(n9644), .op(n9645) );
  mux2_1 U10903 ( .ip1(\cache_data_A[3][83] ), .ip2(n9789), .s(n9645), .op(
        n6917) );
  mux2_1 U10904 ( .ip1(\cache_data_A[3][84] ), .ip2(n9790), .s(n9645), .op(
        n6916) );
  mux2_1 U10905 ( .ip1(\cache_data_A[3][85] ), .ip2(n9791), .s(n9645), .op(
        n6915) );
  mux2_1 U10906 ( .ip1(\cache_data_A[3][86] ), .ip2(n9792), .s(n9645), .op(
        n6914) );
  mux2_1 U10907 ( .ip1(\cache_data_A[3][87] ), .ip2(n9794), .s(n9645), .op(
        n6913) );
  mux2_1 U10908 ( .ip1(\cache_data_A[3][88] ), .ip2(n9795), .s(n9644), .op(
        n6912) );
  mux2_1 U10909 ( .ip1(\cache_data_A[3][89] ), .ip2(n9796), .s(n9644), .op(
        n6911) );
  mux2_1 U10910 ( .ip1(\cache_data_A[3][90] ), .ip2(n9797), .s(n9645), .op(
        n6910) );
  mux2_1 U10911 ( .ip1(\cache_data_A[3][91] ), .ip2(n9798), .s(n9645), .op(
        n6909) );
  mux2_1 U10912 ( .ip1(\cache_data_A[3][92] ), .ip2(n9799), .s(n9645), .op(
        n6908) );
  mux2_1 U10913 ( .ip1(\cache_data_A[3][93] ), .ip2(n9800), .s(n9645), .op(
        n6907) );
  mux2_1 U10914 ( .ip1(\cache_data_A[3][94] ), .ip2(n9801), .s(n9645), .op(
        n6906) );
  mux2_1 U10915 ( .ip1(\cache_data_A[3][95] ), .ip2(n9803), .s(n9645), .op(
        n6905) );
  nor2_1 U10916 ( .ip1(n9866), .ip2(n9672), .op(n9646) );
  mux2_1 U10917 ( .ip1(\cache_data_A[3][96] ), .ip2(n9770), .s(n9646), .op(
        n6904) );
  mux2_1 U10918 ( .ip1(\cache_data_A[3][97] ), .ip2(n9771), .s(n9646), .op(
        n6903) );
  mux2_1 U10919 ( .ip1(\cache_data_A[3][98] ), .ip2(n9772), .s(n9646), .op(
        n6902) );
  mux2_1 U10920 ( .ip1(\cache_data_A[3][99] ), .ip2(n9773), .s(n9646), .op(
        n6901) );
  mux2_1 U10921 ( .ip1(\cache_data_A[3][100] ), .ip2(n9774), .s(n9646), .op(
        n6900) );
  mux2_1 U10922 ( .ip1(\cache_data_A[3][101] ), .ip2(n9775), .s(n9646), .op(
        n6899) );
  mux2_1 U10923 ( .ip1(\cache_data_A[3][102] ), .ip2(n9776), .s(n9646), .op(
        n6898) );
  mux2_1 U10924 ( .ip1(\cache_data_A[3][103] ), .ip2(n9777), .s(n9646), .op(
        n6897) );
  mux2_1 U10925 ( .ip1(\cache_data_A[3][104] ), .ip2(n9778), .s(n9646), .op(
        n6896) );
  mux2_1 U10926 ( .ip1(\cache_data_A[3][105] ), .ip2(n9779), .s(n9646), .op(
        n6895) );
  mux2_1 U10927 ( .ip1(\cache_data_A[3][106] ), .ip2(n9780), .s(n9646), .op(
        n6894) );
  mux2_1 U10928 ( .ip1(\cache_data_A[3][107] ), .ip2(n9781), .s(n9646), .op(
        n6893) );
  mux2_1 U10929 ( .ip1(\cache_data_A[3][108] ), .ip2(n9782), .s(n9646), .op(
        n6892) );
  mux2_1 U10930 ( .ip1(\cache_data_A[3][109] ), .ip2(n9783), .s(n9646), .op(
        n6891) );
  mux2_1 U10931 ( .ip1(\cache_data_A[3][110] ), .ip2(n9784), .s(n9646), .op(
        n6890) );
  mux2_1 U10932 ( .ip1(\cache_data_A[3][111] ), .ip2(n9785), .s(n9646), .op(
        n6889) );
  mux2_1 U10933 ( .ip1(\cache_data_A[3][112] ), .ip2(n9786), .s(n9646), .op(
        n6888) );
  mux2_1 U10934 ( .ip1(\cache_data_A[3][113] ), .ip2(n9787), .s(n9646), .op(
        n6887) );
  mux2_1 U10935 ( .ip1(\cache_data_A[3][114] ), .ip2(n9788), .s(n9646), .op(
        n6886) );
  buf_1 U10936 ( .ip(n9646), .op(n9647) );
  mux2_1 U10937 ( .ip1(\cache_data_A[3][115] ), .ip2(n9789), .s(n9647), .op(
        n6885) );
  mux2_1 U10938 ( .ip1(\cache_data_A[3][116] ), .ip2(n9790), .s(n9647), .op(
        n6884) );
  mux2_1 U10939 ( .ip1(\cache_data_A[3][117] ), .ip2(n9791), .s(n9647), .op(
        n6883) );
  mux2_1 U10940 ( .ip1(\cache_data_A[3][118] ), .ip2(n9792), .s(n9647), .op(
        n6882) );
  mux2_1 U10941 ( .ip1(\cache_data_A[3][119] ), .ip2(n9794), .s(n9647), .op(
        n6881) );
  mux2_1 U10942 ( .ip1(\cache_data_A[3][120] ), .ip2(n9795), .s(n9646), .op(
        n6880) );
  mux2_1 U10943 ( .ip1(\cache_data_A[3][121] ), .ip2(n9796), .s(n9646), .op(
        n6879) );
  mux2_1 U10944 ( .ip1(\cache_data_A[3][122] ), .ip2(n9797), .s(n9647), .op(
        n6878) );
  mux2_1 U10945 ( .ip1(\cache_data_A[3][123] ), .ip2(n9798), .s(n9647), .op(
        n6877) );
  mux2_1 U10946 ( .ip1(\cache_data_A[3][124] ), .ip2(n9799), .s(n9647), .op(
        n6876) );
  mux2_1 U10947 ( .ip1(\cache_data_A[3][125] ), .ip2(n9800), .s(n9647), .op(
        n6875) );
  mux2_1 U10948 ( .ip1(\cache_data_A[3][126] ), .ip2(n9801), .s(n9647), .op(
        n6874) );
  mux2_1 U10949 ( .ip1(\cache_data_A[3][127] ), .ip2(n9803), .s(n9647), .op(
        n6873) );
  nand2_1 U10950 ( .ip1(n9744), .ip2(n9675), .op(n9648) );
  mux2_1 U10951 ( .ip1(n9778), .ip2(\cache_data_A[4][8] ), .s(n9648), .op(
        n6872) );
  mux2_1 U10952 ( .ip1(n9779), .ip2(\cache_data_A[4][9] ), .s(n9648), .op(
        n6871) );
  mux2_1 U10953 ( .ip1(n9780), .ip2(\cache_data_A[4][10] ), .s(n9648), .op(
        n6870) );
  mux2_1 U10954 ( .ip1(n9781), .ip2(\cache_data_A[4][11] ), .s(n9648), .op(
        n6869) );
  mux2_1 U10955 ( .ip1(n9782), .ip2(\cache_data_A[4][12] ), .s(n9648), .op(
        n6868) );
  mux2_1 U10956 ( .ip1(n9783), .ip2(\cache_data_A[4][13] ), .s(n9648), .op(
        n6867) );
  mux2_1 U10957 ( .ip1(n9784), .ip2(\cache_data_A[4][14] ), .s(n9648), .op(
        n6866) );
  mux2_1 U10958 ( .ip1(n9785), .ip2(\cache_data_A[4][15] ), .s(n9648), .op(
        n6865) );
  mux2_1 U10959 ( .ip1(n9786), .ip2(\cache_data_A[4][16] ), .s(n9648), .op(
        n6864) );
  mux2_1 U10960 ( .ip1(n9787), .ip2(\cache_data_A[4][17] ), .s(n9648), .op(
        n6863) );
  mux2_1 U10961 ( .ip1(n9788), .ip2(\cache_data_A[4][18] ), .s(n9648), .op(
        n6862) );
  mux2_1 U10962 ( .ip1(n9789), .ip2(\cache_data_A[4][19] ), .s(n9648), .op(
        n6861) );
  mux2_1 U10963 ( .ip1(n9790), .ip2(\cache_data_A[4][20] ), .s(n9648), .op(
        n6860) );
  mux2_1 U10964 ( .ip1(n9791), .ip2(\cache_data_A[4][21] ), .s(n9648), .op(
        n6859) );
  mux2_1 U10965 ( .ip1(n9792), .ip2(\cache_data_A[4][22] ), .s(n9648), .op(
        n6858) );
  mux2_1 U10966 ( .ip1(n9794), .ip2(\cache_data_A[4][23] ), .s(n9648), .op(
        n6857) );
  mux2_1 U10967 ( .ip1(n9795), .ip2(\cache_data_A[4][24] ), .s(n9648), .op(
        n6856) );
  mux2_1 U10968 ( .ip1(n9796), .ip2(\cache_data_A[4][25] ), .s(n9648), .op(
        n6855) );
  mux2_1 U10969 ( .ip1(n9797), .ip2(\cache_data_A[4][26] ), .s(n9648), .op(
        n6854) );
  buf_1 U10970 ( .ip(n9648), .op(n9649) );
  mux2_1 U10971 ( .ip1(n9798), .ip2(\cache_data_A[4][27] ), .s(n9649), .op(
        n6853) );
  mux2_1 U10972 ( .ip1(n9799), .ip2(\cache_data_A[4][28] ), .s(n9649), .op(
        n6852) );
  mux2_1 U10973 ( .ip1(n9800), .ip2(\cache_data_A[4][29] ), .s(n9649), .op(
        n6851) );
  mux2_1 U10974 ( .ip1(n9801), .ip2(\cache_data_A[4][30] ), .s(n9649), .op(
        n6850) );
  mux2_1 U10975 ( .ip1(n9803), .ip2(\cache_data_A[4][31] ), .s(n9649), .op(
        n6849) );
  mux2_1 U10976 ( .ip1(n9770), .ip2(\cache_data_A[4][0] ), .s(n9648), .op(
        n6848) );
  mux2_1 U10977 ( .ip1(n9771), .ip2(\cache_data_A[4][1] ), .s(n9648), .op(
        n6847) );
  mux2_1 U10978 ( .ip1(n9772), .ip2(\cache_data_A[4][2] ), .s(n9649), .op(
        n6846) );
  mux2_1 U10979 ( .ip1(n9773), .ip2(\cache_data_A[4][3] ), .s(n9649), .op(
        n6845) );
  mux2_1 U10980 ( .ip1(n9774), .ip2(\cache_data_A[4][4] ), .s(n9649), .op(
        n6844) );
  mux2_1 U10981 ( .ip1(n9775), .ip2(\cache_data_A[4][5] ), .s(n9649), .op(
        n6843) );
  mux2_1 U10982 ( .ip1(n9776), .ip2(\cache_data_A[4][6] ), .s(n9649), .op(
        n6842) );
  mux2_1 U10983 ( .ip1(n9777), .ip2(\cache_data_A[4][7] ), .s(n9649), .op(
        n6841) );
  nand2_1 U10984 ( .ip1(n9744), .ip2(n9678), .op(n9650) );
  mux2_1 U10985 ( .ip1(n9812), .ip2(\cache_data_A[4][32] ), .s(n9650), .op(
        n6840) );
  mux2_1 U10986 ( .ip1(n9813), .ip2(\cache_data_A[4][33] ), .s(n9650), .op(
        n6839) );
  mux2_1 U10987 ( .ip1(n9814), .ip2(\cache_data_A[4][34] ), .s(n9650), .op(
        n6838) );
  mux2_1 U10988 ( .ip1(n9815), .ip2(\cache_data_A[4][35] ), .s(n9650), .op(
        n6837) );
  mux2_1 U10989 ( .ip1(n9816), .ip2(\cache_data_A[4][36] ), .s(n9650), .op(
        n6836) );
  mux2_1 U10990 ( .ip1(n9817), .ip2(\cache_data_A[4][37] ), .s(n9650), .op(
        n6835) );
  mux2_1 U10991 ( .ip1(n9818), .ip2(\cache_data_A[4][38] ), .s(n9650), .op(
        n6834) );
  mux2_1 U10992 ( .ip1(n9819), .ip2(\cache_data_A[4][39] ), .s(n9650), .op(
        n6833) );
  mux2_1 U10993 ( .ip1(n9820), .ip2(\cache_data_A[4][40] ), .s(n9650), .op(
        n6832) );
  mux2_1 U10994 ( .ip1(n9821), .ip2(\cache_data_A[4][41] ), .s(n9650), .op(
        n6831) );
  buf_1 U10995 ( .ip(n9650), .op(n9651) );
  mux2_1 U10996 ( .ip1(n9822), .ip2(\cache_data_A[4][42] ), .s(n9651), .op(
        n6830) );
  mux2_1 U10997 ( .ip1(n9823), .ip2(\cache_data_A[4][43] ), .s(n9650), .op(
        n6829) );
  mux2_1 U10998 ( .ip1(n9824), .ip2(\cache_data_A[4][44] ), .s(n9650), .op(
        n6828) );
  mux2_1 U10999 ( .ip1(n9825), .ip2(\cache_data_A[4][45] ), .s(n9650), .op(
        n6827) );
  mux2_1 U11000 ( .ip1(n9826), .ip2(\cache_data_A[4][46] ), .s(n9650), .op(
        n6826) );
  mux2_1 U11001 ( .ip1(n9827), .ip2(\cache_data_A[4][47] ), .s(n9650), .op(
        n6825) );
  mux2_1 U11002 ( .ip1(n9828), .ip2(\cache_data_A[4][48] ), .s(n9651), .op(
        n6824) );
  mux2_1 U11003 ( .ip1(n9829), .ip2(\cache_data_A[4][49] ), .s(n9651), .op(
        n6823) );
  mux2_1 U11004 ( .ip1(n9830), .ip2(\cache_data_A[4][50] ), .s(n9651), .op(
        n6822) );
  mux2_1 U11005 ( .ip1(n9831), .ip2(\cache_data_A[4][51] ), .s(n9650), .op(
        n6821) );
  mux2_1 U11006 ( .ip1(n9832), .ip2(\cache_data_A[4][52] ), .s(n9650), .op(
        n6820) );
  mux2_1 U11007 ( .ip1(n9833), .ip2(\cache_data_A[4][53] ), .s(n9650), .op(
        n6819) );
  mux2_1 U11008 ( .ip1(n9835), .ip2(\cache_data_A[4][54] ), .s(n9650), .op(
        n6818) );
  mux2_1 U11009 ( .ip1(n9836), .ip2(\cache_data_A[4][55] ), .s(n9650), .op(
        n6817) );
  mux2_1 U11010 ( .ip1(n9837), .ip2(\cache_data_A[4][56] ), .s(n9650), .op(
        n6816) );
  mux2_1 U11011 ( .ip1(n9838), .ip2(\cache_data_A[4][57] ), .s(n9651), .op(
        n6815) );
  mux2_1 U11012 ( .ip1(n9839), .ip2(\cache_data_A[4][58] ), .s(n9651), .op(
        n6814) );
  mux2_1 U11013 ( .ip1(n9840), .ip2(\cache_data_A[4][59] ), .s(n9651), .op(
        n6813) );
  mux2_1 U11014 ( .ip1(n9841), .ip2(\cache_data_A[4][60] ), .s(n9651), .op(
        n6812) );
  mux2_1 U11015 ( .ip1(n9842), .ip2(\cache_data_A[4][61] ), .s(n9651), .op(
        n6811) );
  mux2_1 U11016 ( .ip1(n9843), .ip2(\cache_data_A[4][62] ), .s(n9651), .op(
        n6810) );
  mux2_1 U11017 ( .ip1(n9845), .ip2(\cache_data_A[4][63] ), .s(n9651), .op(
        n6809) );
  nor2_1 U11018 ( .ip1(n9868), .ip2(n9681), .op(n9652) );
  mux2_1 U11019 ( .ip1(\cache_data_A[4][64] ), .ip2(n9770), .s(n9652), .op(
        n6808) );
  mux2_1 U11020 ( .ip1(\cache_data_A[4][65] ), .ip2(n9813), .s(n9652), .op(
        n6807) );
  mux2_1 U11021 ( .ip1(\cache_data_A[4][66] ), .ip2(n9814), .s(n9652), .op(
        n6806) );
  mux2_1 U11022 ( .ip1(\cache_data_A[4][67] ), .ip2(n9815), .s(n9652), .op(
        n6805) );
  mux2_1 U11023 ( .ip1(\cache_data_A[4][68] ), .ip2(n9816), .s(n9652), .op(
        n6804) );
  mux2_1 U11024 ( .ip1(\cache_data_A[4][69] ), .ip2(n9817), .s(n9652), .op(
        n6803) );
  mux2_1 U11025 ( .ip1(\cache_data_A[4][70] ), .ip2(n9818), .s(n9652), .op(
        n6802) );
  mux2_1 U11026 ( .ip1(\cache_data_A[4][71] ), .ip2(n9819), .s(n9652), .op(
        n6801) );
  mux2_1 U11027 ( .ip1(\cache_data_A[4][72] ), .ip2(n9820), .s(n9652), .op(
        n6800) );
  buf_1 U11028 ( .ip(n9652), .op(n9653) );
  mux2_1 U11029 ( .ip1(\cache_data_A[4][73] ), .ip2(n9821), .s(n9653), .op(
        n6799) );
  mux2_1 U11030 ( .ip1(\cache_data_A[4][74] ), .ip2(n9822), .s(n9653), .op(
        n6798) );
  mux2_1 U11031 ( .ip1(\cache_data_A[4][75] ), .ip2(n9823), .s(n9652), .op(
        n6797) );
  mux2_1 U11032 ( .ip1(\cache_data_A[4][76] ), .ip2(n9824), .s(n9652), .op(
        n6796) );
  mux2_1 U11033 ( .ip1(\cache_data_A[4][77] ), .ip2(n9825), .s(n9653), .op(
        n6795) );
  mux2_1 U11034 ( .ip1(\cache_data_A[4][78] ), .ip2(n9826), .s(n9652), .op(
        n6794) );
  mux2_1 U11035 ( .ip1(\cache_data_A[4][79] ), .ip2(n9827), .s(n9652), .op(
        n6793) );
  mux2_1 U11036 ( .ip1(\cache_data_A[4][80] ), .ip2(n9828), .s(n9652), .op(
        n6792) );
  mux2_1 U11037 ( .ip1(\cache_data_A[4][81] ), .ip2(n9787), .s(n9652), .op(
        n6791) );
  mux2_1 U11038 ( .ip1(\cache_data_A[4][82] ), .ip2(n9788), .s(n9652), .op(
        n6790) );
  mux2_1 U11039 ( .ip1(\cache_data_A[4][83] ), .ip2(n9831), .s(n9652), .op(
        n6789) );
  mux2_1 U11040 ( .ip1(\cache_data_A[4][84] ), .ip2(n9832), .s(n9652), .op(
        n6788) );
  mux2_1 U11041 ( .ip1(\cache_data_A[4][85] ), .ip2(n9833), .s(n9652), .op(
        n6787) );
  mux2_1 U11042 ( .ip1(\cache_data_A[4][86] ), .ip2(n9835), .s(n9652), .op(
        n6786) );
  mux2_1 U11043 ( .ip1(\cache_data_A[4][87] ), .ip2(n9836), .s(n9652), .op(
        n6785) );
  mux2_1 U11044 ( .ip1(\cache_data_A[4][88] ), .ip2(n9837), .s(n9653), .op(
        n6784) );
  mux2_1 U11045 ( .ip1(\cache_data_A[4][89] ), .ip2(n9796), .s(n9653), .op(
        n6783) );
  mux2_1 U11046 ( .ip1(\cache_data_A[4][90] ), .ip2(n9797), .s(n9653), .op(
        n6782) );
  mux2_1 U11047 ( .ip1(\cache_data_A[4][91] ), .ip2(n9798), .s(n9653), .op(
        n6781) );
  mux2_1 U11048 ( .ip1(\cache_data_A[4][92] ), .ip2(n9799), .s(n9653), .op(
        n6780) );
  mux2_1 U11049 ( .ip1(\cache_data_A[4][93] ), .ip2(n9800), .s(n9653), .op(
        n6779) );
  mux2_1 U11050 ( .ip1(\cache_data_A[4][94] ), .ip2(n9801), .s(n9653), .op(
        n6778) );
  mux2_1 U11051 ( .ip1(\cache_data_A[4][95] ), .ip2(n9803), .s(n9653), .op(
        n6777) );
  nand2_1 U11052 ( .ip1(n9744), .ip2(n9684), .op(n9654) );
  mux2_1 U11053 ( .ip1(n9823), .ip2(\cache_data_A[4][107] ), .s(n9654), .op(
        n6776) );
  mux2_1 U11054 ( .ip1(n9824), .ip2(\cache_data_A[4][108] ), .s(n9654), .op(
        n6775) );
  mux2_1 U11055 ( .ip1(n9825), .ip2(\cache_data_A[4][109] ), .s(n9654), .op(
        n6774) );
  mux2_1 U11056 ( .ip1(n9826), .ip2(\cache_data_A[4][110] ), .s(n9654), .op(
        n6773) );
  mux2_1 U11057 ( .ip1(n9827), .ip2(\cache_data_A[4][111] ), .s(n9654), .op(
        n6772) );
  mux2_1 U11058 ( .ip1(n9828), .ip2(\cache_data_A[4][112] ), .s(n9654), .op(
        n6771) );
  mux2_1 U11059 ( .ip1(n9829), .ip2(\cache_data_A[4][113] ), .s(n9654), .op(
        n6770) );
  mux2_1 U11060 ( .ip1(n9830), .ip2(\cache_data_A[4][114] ), .s(n9654), .op(
        n6769) );
  mux2_1 U11061 ( .ip1(n9831), .ip2(\cache_data_A[4][115] ), .s(n9654), .op(
        n6768) );
  mux2_1 U11062 ( .ip1(n9832), .ip2(\cache_data_A[4][116] ), .s(n9654), .op(
        n6767) );
  mux2_1 U11063 ( .ip1(n9833), .ip2(\cache_data_A[4][117] ), .s(n9654), .op(
        n6766) );
  mux2_1 U11064 ( .ip1(n9835), .ip2(\cache_data_A[4][118] ), .s(n9654), .op(
        n6765) );
  mux2_1 U11065 ( .ip1(n9836), .ip2(\cache_data_A[4][119] ), .s(n9654), .op(
        n6764) );
  mux2_1 U11066 ( .ip1(n9837), .ip2(\cache_data_A[4][120] ), .s(n9654), .op(
        n6763) );
  mux2_1 U11067 ( .ip1(n9838), .ip2(\cache_data_A[4][121] ), .s(n9654), .op(
        n6762) );
  mux2_1 U11068 ( .ip1(n9839), .ip2(\cache_data_A[4][122] ), .s(n9654), .op(
        n6761) );
  mux2_1 U11069 ( .ip1(n9840), .ip2(\cache_data_A[4][123] ), .s(n9654), .op(
        n6760) );
  mux2_1 U11070 ( .ip1(n9841), .ip2(\cache_data_A[4][124] ), .s(n9654), .op(
        n6759) );
  mux2_1 U11071 ( .ip1(n9842), .ip2(\cache_data_A[4][125] ), .s(n9654), .op(
        n6758) );
  buf_1 U11072 ( .ip(n9654), .op(n9655) );
  mux2_1 U11073 ( .ip1(n9843), .ip2(\cache_data_A[4][126] ), .s(n9655), .op(
        n6757) );
  mux2_1 U11074 ( .ip1(n9845), .ip2(\cache_data_A[4][127] ), .s(n9655), .op(
        n6756) );
  mux2_1 U11075 ( .ip1(n9812), .ip2(\cache_data_A[4][96] ), .s(n9655), .op(
        n6755) );
  mux2_1 U11076 ( .ip1(n9813), .ip2(\cache_data_A[4][97] ), .s(n9655), .op(
        n6754) );
  mux2_1 U11077 ( .ip1(n9814), .ip2(\cache_data_A[4][98] ), .s(n9655), .op(
        n6753) );
  mux2_1 U11078 ( .ip1(n9815), .ip2(\cache_data_A[4][99] ), .s(n9654), .op(
        n6752) );
  mux2_1 U11079 ( .ip1(n9816), .ip2(\cache_data_A[4][100] ), .s(n9654), .op(
        n6751) );
  mux2_1 U11080 ( .ip1(n9817), .ip2(\cache_data_A[4][101] ), .s(n9655), .op(
        n6750) );
  mux2_1 U11081 ( .ip1(n9818), .ip2(\cache_data_A[4][102] ), .s(n9655), .op(
        n6749) );
  mux2_1 U11082 ( .ip1(n9819), .ip2(\cache_data_A[4][103] ), .s(n9655), .op(
        n6748) );
  mux2_1 U11083 ( .ip1(n9820), .ip2(\cache_data_A[4][104] ), .s(n9655), .op(
        n6747) );
  mux2_1 U11084 ( .ip1(n9821), .ip2(\cache_data_A[4][105] ), .s(n9655), .op(
        n6746) );
  mux2_1 U11085 ( .ip1(n9822), .ip2(\cache_data_A[4][106] ), .s(n9655), .op(
        n6745) );
  nor2_1 U11086 ( .ip1(n9870), .ip2(n9665), .op(n9656) );
  mux2_1 U11087 ( .ip1(\cache_data_A[5][0] ), .ip2(n9812), .s(n9656), .op(
        n6744) );
  mux2_1 U11088 ( .ip1(\cache_data_A[5][1] ), .ip2(n9771), .s(n9656), .op(
        n6743) );
  mux2_1 U11089 ( .ip1(\cache_data_A[5][2] ), .ip2(n9772), .s(n9656), .op(
        n6742) );
  mux2_1 U11090 ( .ip1(\cache_data_A[5][3] ), .ip2(n9773), .s(n9656), .op(
        n6741) );
  mux2_1 U11091 ( .ip1(\cache_data_A[5][4] ), .ip2(n9774), .s(n9656), .op(
        n6740) );
  mux2_1 U11092 ( .ip1(\cache_data_A[5][5] ), .ip2(n9775), .s(n9656), .op(
        n6739) );
  mux2_1 U11093 ( .ip1(\cache_data_A[5][6] ), .ip2(n9776), .s(n9656), .op(
        n6738) );
  mux2_1 U11094 ( .ip1(\cache_data_A[5][7] ), .ip2(n9777), .s(n9656), .op(
        n6737) );
  mux2_1 U11095 ( .ip1(\cache_data_A[5][8] ), .ip2(n9778), .s(n9656), .op(
        n6736) );
  mux2_1 U11096 ( .ip1(\cache_data_A[5][9] ), .ip2(n9779), .s(n9656), .op(
        n6735) );
  mux2_1 U11097 ( .ip1(\cache_data_A[5][10] ), .ip2(n9780), .s(n9656), .op(
        n6734) );
  mux2_1 U11098 ( .ip1(\cache_data_A[5][11] ), .ip2(n9781), .s(n9656), .op(
        n6733) );
  mux2_1 U11099 ( .ip1(\cache_data_A[5][12] ), .ip2(n9782), .s(n9656), .op(
        n6732) );
  mux2_1 U11100 ( .ip1(\cache_data_A[5][13] ), .ip2(n9783), .s(n9656), .op(
        n6731) );
  mux2_1 U11101 ( .ip1(\cache_data_A[5][14] ), .ip2(n9784), .s(n9656), .op(
        n6730) );
  mux2_1 U11102 ( .ip1(\cache_data_A[5][15] ), .ip2(n9785), .s(n9656), .op(
        n6729) );
  mux2_1 U11103 ( .ip1(\cache_data_A[5][16] ), .ip2(n9786), .s(n9656), .op(
        n6728) );
  mux2_1 U11104 ( .ip1(\cache_data_A[5][17] ), .ip2(n9829), .s(n9656), .op(
        n6727) );
  mux2_1 U11105 ( .ip1(\cache_data_A[5][18] ), .ip2(n9830), .s(n9656), .op(
        n6726) );
  buf_1 U11106 ( .ip(n9656), .op(n9657) );
  mux2_1 U11107 ( .ip1(\cache_data_A[5][19] ), .ip2(n9831), .s(n9657), .op(
        n6725) );
  mux2_1 U11108 ( .ip1(\cache_data_A[5][20] ), .ip2(n9832), .s(n9657), .op(
        n6724) );
  mux2_1 U11109 ( .ip1(\cache_data_A[5][21] ), .ip2(n9833), .s(n9657), .op(
        n6723) );
  mux2_1 U11110 ( .ip1(\cache_data_A[5][22] ), .ip2(n9835), .s(n9657), .op(
        n6722) );
  mux2_1 U11111 ( .ip1(\cache_data_A[5][23] ), .ip2(n9836), .s(n9657), .op(
        n6721) );
  mux2_1 U11112 ( .ip1(\cache_data_A[5][24] ), .ip2(n9837), .s(n9656), .op(
        n6720) );
  mux2_1 U11113 ( .ip1(\cache_data_A[5][25] ), .ip2(n9838), .s(n9656), .op(
        n6719) );
  mux2_1 U11114 ( .ip1(\cache_data_A[5][26] ), .ip2(n9839), .s(n9657), .op(
        n6718) );
  mux2_1 U11115 ( .ip1(\cache_data_A[5][27] ), .ip2(n9840), .s(n9657), .op(
        n6717) );
  mux2_1 U11116 ( .ip1(\cache_data_A[5][28] ), .ip2(n9841), .s(n9657), .op(
        n6716) );
  mux2_1 U11117 ( .ip1(\cache_data_A[5][29] ), .ip2(n9842), .s(n9657), .op(
        n6715) );
  mux2_1 U11118 ( .ip1(\cache_data_A[5][30] ), .ip2(n9843), .s(n9657), .op(
        n6714) );
  mux2_1 U11119 ( .ip1(\cache_data_A[5][31] ), .ip2(n9845), .s(n9657), .op(
        n6713) );
  nand2_1 U11120 ( .ip1(n9753), .ip2(n9678), .op(n9658) );
  mux2_1 U11121 ( .ip1(n9812), .ip2(\cache_data_A[5][32] ), .s(n9658), .op(
        n6712) );
  mux2_1 U11122 ( .ip1(n9813), .ip2(\cache_data_A[5][33] ), .s(n9658), .op(
        n6711) );
  mux2_1 U11123 ( .ip1(n9814), .ip2(\cache_data_A[5][34] ), .s(n9658), .op(
        n6710) );
  mux2_1 U11124 ( .ip1(n9815), .ip2(\cache_data_A[5][35] ), .s(n9658), .op(
        n6709) );
  mux2_1 U11125 ( .ip1(n9816), .ip2(\cache_data_A[5][36] ), .s(n9658), .op(
        n6708) );
  mux2_1 U11126 ( .ip1(n9817), .ip2(\cache_data_A[5][37] ), .s(n9658), .op(
        n6707) );
  mux2_1 U11127 ( .ip1(n9818), .ip2(\cache_data_A[5][38] ), .s(n9658), .op(
        n6706) );
  mux2_1 U11128 ( .ip1(n9819), .ip2(\cache_data_A[5][39] ), .s(n9658), .op(
        n6705) );
  mux2_1 U11129 ( .ip1(n9820), .ip2(\cache_data_A[5][40] ), .s(n9658), .op(
        n6704) );
  buf_1 U11130 ( .ip(n9658), .op(n9659) );
  mux2_1 U11131 ( .ip1(n9821), .ip2(\cache_data_A[5][41] ), .s(n9659), .op(
        n6703) );
  mux2_1 U11132 ( .ip1(n9822), .ip2(\cache_data_A[5][42] ), .s(n9658), .op(
        n6702) );
  mux2_1 U11133 ( .ip1(n9823), .ip2(\cache_data_A[5][43] ), .s(n9658), .op(
        n6701) );
  mux2_1 U11134 ( .ip1(n9824), .ip2(\cache_data_A[5][44] ), .s(n9658), .op(
        n6700) );
  mux2_1 U11135 ( .ip1(n9825), .ip2(\cache_data_A[5][45] ), .s(n9658), .op(
        n6699) );
  mux2_1 U11136 ( .ip1(n9826), .ip2(\cache_data_A[5][46] ), .s(n9658), .op(
        n6698) );
  mux2_1 U11137 ( .ip1(n9827), .ip2(\cache_data_A[5][47] ), .s(n9658), .op(
        n6697) );
  mux2_1 U11138 ( .ip1(n9828), .ip2(\cache_data_A[5][48] ), .s(n9658), .op(
        n6696) );
  mux2_1 U11139 ( .ip1(n9829), .ip2(\cache_data_A[5][49] ), .s(n9658), .op(
        n6695) );
  mux2_1 U11140 ( .ip1(n9830), .ip2(\cache_data_A[5][50] ), .s(n9658), .op(
        n6694) );
  mux2_1 U11141 ( .ip1(n9831), .ip2(\cache_data_A[5][51] ), .s(n9658), .op(
        n6693) );
  mux2_1 U11142 ( .ip1(n9832), .ip2(\cache_data_A[5][52] ), .s(n9658), .op(
        n6692) );
  mux2_1 U11143 ( .ip1(n9833), .ip2(\cache_data_A[5][53] ), .s(n9658), .op(
        n6691) );
  mux2_1 U11144 ( .ip1(n9835), .ip2(\cache_data_A[5][54] ), .s(n9659), .op(
        n6690) );
  mux2_1 U11145 ( .ip1(n9836), .ip2(\cache_data_A[5][55] ), .s(n9659), .op(
        n6689) );
  mux2_1 U11146 ( .ip1(n9837), .ip2(\cache_data_A[5][56] ), .s(n9659), .op(
        n6688) );
  mux2_1 U11147 ( .ip1(n9838), .ip2(\cache_data_A[5][57] ), .s(n9659), .op(
        n6687) );
  mux2_1 U11148 ( .ip1(n9839), .ip2(\cache_data_A[5][58] ), .s(n9659), .op(
        n6686) );
  mux2_1 U11149 ( .ip1(n9840), .ip2(\cache_data_A[5][59] ), .s(n9659), .op(
        n6685) );
  mux2_1 U11150 ( .ip1(n9841), .ip2(\cache_data_A[5][60] ), .s(n9659), .op(
        n6684) );
  mux2_1 U11151 ( .ip1(n9842), .ip2(\cache_data_A[5][61] ), .s(n9659), .op(
        n6683) );
  mux2_1 U11152 ( .ip1(n9843), .ip2(\cache_data_A[5][62] ), .s(n9659), .op(
        n6682) );
  mux2_1 U11153 ( .ip1(n9845), .ip2(\cache_data_A[5][63] ), .s(n9659), .op(
        n6681) );
  nand2_1 U11154 ( .ip1(n9753), .ip2(n9660), .op(n9661) );
  mux2_1 U11155 ( .ip1(n9826), .ip2(\cache_data_A[5][78] ), .s(n9661), .op(
        n6680) );
  mux2_1 U11156 ( .ip1(n9827), .ip2(\cache_data_A[5][79] ), .s(n9661), .op(
        n6679) );
  mux2_1 U11157 ( .ip1(n9828), .ip2(\cache_data_A[5][80] ), .s(n9661), .op(
        n6678) );
  mux2_1 U11158 ( .ip1(n9829), .ip2(\cache_data_A[5][81] ), .s(n9661), .op(
        n6677) );
  mux2_1 U11159 ( .ip1(n9830), .ip2(\cache_data_A[5][82] ), .s(n9661), .op(
        n6676) );
  mux2_1 U11160 ( .ip1(n9789), .ip2(\cache_data_A[5][83] ), .s(n9661), .op(
        n6675) );
  mux2_1 U11161 ( .ip1(n9832), .ip2(\cache_data_A[5][84] ), .s(n9661), .op(
        n6674) );
  mux2_1 U11162 ( .ip1(n9833), .ip2(\cache_data_A[5][85] ), .s(n9661), .op(
        n6673) );
  mux2_1 U11163 ( .ip1(n9835), .ip2(\cache_data_A[5][86] ), .s(n9661), .op(
        n6672) );
  buf_1 U11164 ( .ip(n9661), .op(n9662) );
  mux2_1 U11165 ( .ip1(n9836), .ip2(\cache_data_A[5][87] ), .s(n9662), .op(
        n6671) );
  mux2_1 U11166 ( .ip1(n9837), .ip2(\cache_data_A[5][88] ), .s(n9661), .op(
        n6670) );
  mux2_1 U11167 ( .ip1(n9838), .ip2(\cache_data_A[5][89] ), .s(n9661), .op(
        n6669) );
  mux2_1 U11168 ( .ip1(n9839), .ip2(\cache_data_A[5][90] ), .s(n9661), .op(
        n6668) );
  mux2_1 U11169 ( .ip1(n9840), .ip2(\cache_data_A[5][91] ), .s(n9661), .op(
        n6667) );
  mux2_1 U11170 ( .ip1(n9841), .ip2(\cache_data_A[5][92] ), .s(n9661), .op(
        n6666) );
  mux2_1 U11171 ( .ip1(n9842), .ip2(\cache_data_A[5][93] ), .s(n9661), .op(
        n6665) );
  mux2_1 U11172 ( .ip1(n9843), .ip2(\cache_data_A[5][94] ), .s(n9661), .op(
        n6664) );
  mux2_1 U11173 ( .ip1(n9845), .ip2(\cache_data_A[5][95] ), .s(n9661), .op(
        n6663) );
  mux2_1 U11174 ( .ip1(n9812), .ip2(\cache_data_A[5][64] ), .s(n9661), .op(
        n6662) );
  mux2_1 U11175 ( .ip1(n9813), .ip2(\cache_data_A[5][65] ), .s(n9661), .op(
        n6661) );
  mux2_1 U11176 ( .ip1(n9814), .ip2(\cache_data_A[5][66] ), .s(n9661), .op(
        n6660) );
  mux2_1 U11177 ( .ip1(n9815), .ip2(\cache_data_A[5][67] ), .s(n9661), .op(
        n6659) );
  mux2_1 U11178 ( .ip1(n9816), .ip2(\cache_data_A[5][68] ), .s(n9662), .op(
        n6658) );
  mux2_1 U11179 ( .ip1(n9817), .ip2(\cache_data_A[5][69] ), .s(n9662), .op(
        n6657) );
  mux2_1 U11180 ( .ip1(n9818), .ip2(\cache_data_A[5][70] ), .s(n9662), .op(
        n6656) );
  mux2_1 U11181 ( .ip1(n9819), .ip2(\cache_data_A[5][71] ), .s(n9662), .op(
        n6655) );
  mux2_1 U11182 ( .ip1(n9820), .ip2(\cache_data_A[5][72] ), .s(n9662), .op(
        n6654) );
  mux2_1 U11183 ( .ip1(n9821), .ip2(\cache_data_A[5][73] ), .s(n9662), .op(
        n6653) );
  mux2_1 U11184 ( .ip1(n9822), .ip2(\cache_data_A[5][74] ), .s(n9662), .op(
        n6652) );
  mux2_1 U11185 ( .ip1(n9823), .ip2(\cache_data_A[5][75] ), .s(n9662), .op(
        n6651) );
  mux2_1 U11186 ( .ip1(n9824), .ip2(\cache_data_A[5][76] ), .s(n9662), .op(
        n6650) );
  mux2_1 U11187 ( .ip1(n9825), .ip2(\cache_data_A[5][77] ), .s(n9662), .op(
        n6649) );
  nor2_1 U11188 ( .ip1(n9870), .ip2(n9672), .op(n9663) );
  mux2_1 U11189 ( .ip1(\cache_data_A[5][96] ), .ip2(n9770), .s(n9663), .op(
        n6648) );
  mux2_1 U11190 ( .ip1(\cache_data_A[5][97] ), .ip2(n9771), .s(n9663), .op(
        n6647) );
  mux2_1 U11191 ( .ip1(\cache_data_A[5][98] ), .ip2(n9772), .s(n9663), .op(
        n6646) );
  mux2_1 U11192 ( .ip1(\cache_data_A[5][99] ), .ip2(n9773), .s(n9663), .op(
        n6645) );
  mux2_1 U11193 ( .ip1(\cache_data_A[5][100] ), .ip2(n9774), .s(n9663), .op(
        n6644) );
  mux2_1 U11194 ( .ip1(\cache_data_A[5][101] ), .ip2(n9775), .s(n9663), .op(
        n6643) );
  mux2_1 U11195 ( .ip1(\cache_data_A[5][102] ), .ip2(n9776), .s(n9663), .op(
        n6642) );
  mux2_1 U11196 ( .ip1(\cache_data_A[5][103] ), .ip2(n9777), .s(n9663), .op(
        n6641) );
  mux2_1 U11197 ( .ip1(\cache_data_A[5][104] ), .ip2(n9778), .s(n9663), .op(
        n6640) );
  mux2_1 U11198 ( .ip1(\cache_data_A[5][105] ), .ip2(n9779), .s(n9663), .op(
        n6639) );
  mux2_1 U11199 ( .ip1(\cache_data_A[5][106] ), .ip2(n9780), .s(n9663), .op(
        n6638) );
  mux2_1 U11200 ( .ip1(\cache_data_A[5][107] ), .ip2(n9781), .s(n9663), .op(
        n6637) );
  mux2_1 U11201 ( .ip1(\cache_data_A[5][108] ), .ip2(n9782), .s(n9663), .op(
        n6636) );
  mux2_1 U11202 ( .ip1(\cache_data_A[5][109] ), .ip2(n9783), .s(n9663), .op(
        n6635) );
  mux2_1 U11203 ( .ip1(\cache_data_A[5][110] ), .ip2(n9784), .s(n9663), .op(
        n6634) );
  mux2_1 U11204 ( .ip1(\cache_data_A[5][111] ), .ip2(n9785), .s(n9663), .op(
        n6633) );
  mux2_1 U11205 ( .ip1(\cache_data_A[5][112] ), .ip2(n9786), .s(n9663), .op(
        n6632) );
  mux2_1 U11206 ( .ip1(\cache_data_A[5][113] ), .ip2(n9787), .s(n9663), .op(
        n6631) );
  mux2_1 U11207 ( .ip1(\cache_data_A[5][114] ), .ip2(n9788), .s(n9663), .op(
        n6630) );
  buf_1 U11208 ( .ip(n9663), .op(n9664) );
  mux2_1 U11209 ( .ip1(\cache_data_A[5][115] ), .ip2(n9789), .s(n9664), .op(
        n6629) );
  mux2_1 U11210 ( .ip1(\cache_data_A[5][116] ), .ip2(n9790), .s(n9664), .op(
        n6628) );
  mux2_1 U11211 ( .ip1(\cache_data_A[5][117] ), .ip2(n9791), .s(n9664), .op(
        n6627) );
  mux2_1 U11212 ( .ip1(\cache_data_A[5][118] ), .ip2(n9792), .s(n9664), .op(
        n6626) );
  mux2_1 U11213 ( .ip1(\cache_data_A[5][119] ), .ip2(n9794), .s(n9664), .op(
        n6625) );
  mux2_1 U11214 ( .ip1(\cache_data_A[5][120] ), .ip2(n9795), .s(n9663), .op(
        n6624) );
  mux2_1 U11215 ( .ip1(\cache_data_A[5][121] ), .ip2(n9796), .s(n9663), .op(
        n6623) );
  mux2_1 U11216 ( .ip1(\cache_data_A[5][122] ), .ip2(n9797), .s(n9664), .op(
        n6622) );
  mux2_1 U11217 ( .ip1(\cache_data_A[5][123] ), .ip2(n9798), .s(n9664), .op(
        n6621) );
  mux2_1 U11218 ( .ip1(\cache_data_A[5][124] ), .ip2(n9799), .s(n9664), .op(
        n6620) );
  mux2_1 U11219 ( .ip1(\cache_data_A[5][125] ), .ip2(n9800), .s(n9664), .op(
        n6619) );
  mux2_1 U11220 ( .ip1(\cache_data_A[5][126] ), .ip2(n9801), .s(n9664), .op(
        n6618) );
  mux2_1 U11221 ( .ip1(\cache_data_A[5][127] ), .ip2(n9803), .s(n9664), .op(
        n6617) );
  nor2_1 U11222 ( .ip1(n9762), .ip2(n9665), .op(n9666) );
  mux2_1 U11223 ( .ip1(\cache_data_A[6][0] ), .ip2(n9770), .s(n9666), .op(
        n6616) );
  mux2_1 U11224 ( .ip1(\cache_data_A[6][1] ), .ip2(n9771), .s(n9666), .op(
        n6615) );
  mux2_1 U11225 ( .ip1(\cache_data_A[6][2] ), .ip2(n9772), .s(n9666), .op(
        n6614) );
  mux2_1 U11226 ( .ip1(\cache_data_A[6][3] ), .ip2(n9773), .s(n9666), .op(
        n6613) );
  mux2_1 U11227 ( .ip1(\cache_data_A[6][4] ), .ip2(n9774), .s(n9666), .op(
        n6612) );
  mux2_1 U11228 ( .ip1(\cache_data_A[6][5] ), .ip2(n9775), .s(n9666), .op(
        n6611) );
  mux2_1 U11229 ( .ip1(\cache_data_A[6][6] ), .ip2(n9776), .s(n9666), .op(
        n6610) );
  mux2_1 U11230 ( .ip1(\cache_data_A[6][7] ), .ip2(n9777), .s(n9666), .op(
        n6609) );
  mux2_1 U11231 ( .ip1(\cache_data_A[6][8] ), .ip2(n9778), .s(n9666), .op(
        n6608) );
  buf_1 U11232 ( .ip(n9666), .op(n9667) );
  mux2_1 U11233 ( .ip1(\cache_data_A[6][9] ), .ip2(n9779), .s(n9667), .op(
        n6607) );
  mux2_1 U11234 ( .ip1(\cache_data_A[6][10] ), .ip2(n9780), .s(n9667), .op(
        n6606) );
  mux2_1 U11235 ( .ip1(\cache_data_A[6][11] ), .ip2(n9781), .s(n9666), .op(
        n6605) );
  mux2_1 U11236 ( .ip1(\cache_data_A[6][12] ), .ip2(n9782), .s(n9666), .op(
        n6604) );
  mux2_1 U11237 ( .ip1(\cache_data_A[6][13] ), .ip2(n9783), .s(n9667), .op(
        n6603) );
  mux2_1 U11238 ( .ip1(\cache_data_A[6][14] ), .ip2(n9784), .s(n9666), .op(
        n6602) );
  mux2_1 U11239 ( .ip1(\cache_data_A[6][15] ), .ip2(n9785), .s(n9666), .op(
        n6601) );
  mux2_1 U11240 ( .ip1(\cache_data_A[6][16] ), .ip2(n9786), .s(n9666), .op(
        n6600) );
  mux2_1 U11241 ( .ip1(\cache_data_A[6][17] ), .ip2(n9787), .s(n9666), .op(
        n6599) );
  mux2_1 U11242 ( .ip1(\cache_data_A[6][18] ), .ip2(n9788), .s(n9666), .op(
        n6598) );
  mux2_1 U11243 ( .ip1(\cache_data_A[6][19] ), .ip2(n9789), .s(n9666), .op(
        n6597) );
  mux2_1 U11244 ( .ip1(\cache_data_A[6][20] ), .ip2(n9790), .s(n9666), .op(
        n6596) );
  mux2_1 U11245 ( .ip1(\cache_data_A[6][21] ), .ip2(n9791), .s(n9666), .op(
        n6595) );
  mux2_1 U11246 ( .ip1(\cache_data_A[6][22] ), .ip2(n9792), .s(n9666), .op(
        n6594) );
  mux2_1 U11247 ( .ip1(\cache_data_A[6][23] ), .ip2(n9794), .s(n9666), .op(
        n6593) );
  mux2_1 U11248 ( .ip1(\cache_data_A[6][24] ), .ip2(n9795), .s(n9667), .op(
        n6592) );
  mux2_1 U11249 ( .ip1(\cache_data_A[6][25] ), .ip2(n9796), .s(n9667), .op(
        n6591) );
  mux2_1 U11250 ( .ip1(\cache_data_A[6][26] ), .ip2(n9797), .s(n9667), .op(
        n6590) );
  mux2_1 U11251 ( .ip1(\cache_data_A[6][27] ), .ip2(n9798), .s(n9667), .op(
        n6589) );
  mux2_1 U11252 ( .ip1(\cache_data_A[6][28] ), .ip2(n9799), .s(n9667), .op(
        n6588) );
  mux2_1 U11253 ( .ip1(\cache_data_A[6][29] ), .ip2(n9800), .s(n9667), .op(
        n6587) );
  mux2_1 U11254 ( .ip1(\cache_data_A[6][30] ), .ip2(n9801), .s(n9667), .op(
        n6586) );
  mux2_1 U11255 ( .ip1(\cache_data_A[6][31] ), .ip2(n9803), .s(n9667), .op(
        n6585) );
  nand2_1 U11256 ( .ip1(n9765), .ip2(n9678), .op(n9668) );
  mux2_1 U11257 ( .ip1(n9829), .ip2(\cache_data_A[6][49] ), .s(n9668), .op(
        n6584) );
  mux2_1 U11258 ( .ip1(n9830), .ip2(\cache_data_A[6][50] ), .s(n9668), .op(
        n6583) );
  mux2_1 U11259 ( .ip1(n9831), .ip2(\cache_data_A[6][51] ), .s(n9668), .op(
        n6582) );
  mux2_1 U11260 ( .ip1(n9832), .ip2(\cache_data_A[6][52] ), .s(n9668), .op(
        n6581) );
  mux2_1 U11261 ( .ip1(n9833), .ip2(\cache_data_A[6][53] ), .s(n9668), .op(
        n6580) );
  mux2_1 U11262 ( .ip1(n9835), .ip2(\cache_data_A[6][54] ), .s(n9668), .op(
        n6579) );
  mux2_1 U11263 ( .ip1(n9836), .ip2(\cache_data_A[6][55] ), .s(n9668), .op(
        n6578) );
  mux2_1 U11264 ( .ip1(n9837), .ip2(\cache_data_A[6][56] ), .s(n9668), .op(
        n6577) );
  mux2_1 U11265 ( .ip1(n9838), .ip2(\cache_data_A[6][57] ), .s(n9668), .op(
        n6576) );
  mux2_1 U11266 ( .ip1(n9839), .ip2(\cache_data_A[6][58] ), .s(n9668), .op(
        n6575) );
  buf_1 U11267 ( .ip(n9668), .op(n9669) );
  mux2_1 U11268 ( .ip1(n9840), .ip2(\cache_data_A[6][59] ), .s(n9669), .op(
        n6574) );
  mux2_1 U11269 ( .ip1(n9841), .ip2(\cache_data_A[6][60] ), .s(n9668), .op(
        n6573) );
  mux2_1 U11270 ( .ip1(n9842), .ip2(\cache_data_A[6][61] ), .s(n9668), .op(
        n6572) );
  mux2_1 U11271 ( .ip1(n9843), .ip2(\cache_data_A[6][62] ), .s(n9669), .op(
        n6571) );
  mux2_1 U11272 ( .ip1(n9845), .ip2(\cache_data_A[6][63] ), .s(n9668), .op(
        n6570) );
  mux2_1 U11273 ( .ip1(n9812), .ip2(\cache_data_A[6][32] ), .s(n9668), .op(
        n6569) );
  mux2_1 U11274 ( .ip1(n9813), .ip2(\cache_data_A[6][33] ), .s(n9668), .op(
        n6568) );
  mux2_1 U11275 ( .ip1(n9814), .ip2(\cache_data_A[6][34] ), .s(n9668), .op(
        n6567) );
  mux2_1 U11276 ( .ip1(n9815), .ip2(\cache_data_A[6][35] ), .s(n9668), .op(
        n6566) );
  mux2_1 U11277 ( .ip1(n9816), .ip2(\cache_data_A[6][36] ), .s(n9668), .op(
        n6565) );
  mux2_1 U11278 ( .ip1(n9817), .ip2(\cache_data_A[6][37] ), .s(n9668), .op(
        n6564) );
  mux2_1 U11279 ( .ip1(n9818), .ip2(\cache_data_A[6][38] ), .s(n9668), .op(
        n6563) );
  mux2_1 U11280 ( .ip1(n9819), .ip2(\cache_data_A[6][39] ), .s(n9668), .op(
        n6562) );
  mux2_1 U11281 ( .ip1(n9820), .ip2(\cache_data_A[6][40] ), .s(n9669), .op(
        n6561) );
  mux2_1 U11282 ( .ip1(n9821), .ip2(\cache_data_A[6][41] ), .s(n9669), .op(
        n6560) );
  mux2_1 U11283 ( .ip1(n9822), .ip2(\cache_data_A[6][42] ), .s(n9669), .op(
        n6559) );
  mux2_1 U11284 ( .ip1(n9823), .ip2(\cache_data_A[6][43] ), .s(n9669), .op(
        n6558) );
  mux2_1 U11285 ( .ip1(n9824), .ip2(\cache_data_A[6][44] ), .s(n9669), .op(
        n6557) );
  mux2_1 U11286 ( .ip1(n9825), .ip2(\cache_data_A[6][45] ), .s(n9669), .op(
        n6556) );
  mux2_1 U11287 ( .ip1(n9826), .ip2(\cache_data_A[6][46] ), .s(n9669), .op(
        n6555) );
  mux2_1 U11288 ( .ip1(n9827), .ip2(\cache_data_A[6][47] ), .s(n9669), .op(
        n6554) );
  mux2_1 U11289 ( .ip1(n9828), .ip2(\cache_data_A[6][48] ), .s(n9669), .op(
        n6553) );
  nor2_1 U11290 ( .ip1(n9762), .ip2(n9681), .op(n9670) );
  mux2_1 U11291 ( .ip1(\cache_data_A[6][64] ), .ip2(n9770), .s(n9670), .op(
        n6552) );
  mux2_1 U11292 ( .ip1(\cache_data_A[6][65] ), .ip2(n9771), .s(n9670), .op(
        n6551) );
  mux2_1 U11293 ( .ip1(\cache_data_A[6][66] ), .ip2(n9772), .s(n9670), .op(
        n6550) );
  mux2_1 U11294 ( .ip1(\cache_data_A[6][67] ), .ip2(n9773), .s(n9670), .op(
        n6549) );
  mux2_1 U11295 ( .ip1(\cache_data_A[6][68] ), .ip2(n9774), .s(n9670), .op(
        n6548) );
  mux2_1 U11296 ( .ip1(\cache_data_A[6][69] ), .ip2(n9775), .s(n9670), .op(
        n6547) );
  mux2_1 U11297 ( .ip1(\cache_data_A[6][70] ), .ip2(n9776), .s(n9670), .op(
        n6546) );
  mux2_1 U11298 ( .ip1(\cache_data_A[6][71] ), .ip2(n9777), .s(n9670), .op(
        n6545) );
  mux2_1 U11299 ( .ip1(\cache_data_A[6][72] ), .ip2(n9778), .s(n9670), .op(
        n6544) );
  buf_1 U11300 ( .ip(n9670), .op(n9671) );
  mux2_1 U11301 ( .ip1(\cache_data_A[6][73] ), .ip2(n9779), .s(n9671), .op(
        n6543) );
  mux2_1 U11302 ( .ip1(\cache_data_A[6][74] ), .ip2(n9780), .s(n9671), .op(
        n6542) );
  mux2_1 U11303 ( .ip1(\cache_data_A[6][75] ), .ip2(n9781), .s(n9670), .op(
        n6541) );
  mux2_1 U11304 ( .ip1(\cache_data_A[6][76] ), .ip2(n9782), .s(n9670), .op(
        n6540) );
  mux2_1 U11305 ( .ip1(\cache_data_A[6][77] ), .ip2(n9783), .s(n9671), .op(
        n6539) );
  mux2_1 U11306 ( .ip1(\cache_data_A[6][78] ), .ip2(n9784), .s(n9670), .op(
        n6538) );
  mux2_1 U11307 ( .ip1(\cache_data_A[6][79] ), .ip2(n9785), .s(n9670), .op(
        n6537) );
  mux2_1 U11308 ( .ip1(\cache_data_A[6][80] ), .ip2(n9786), .s(n9670), .op(
        n6536) );
  mux2_1 U11309 ( .ip1(\cache_data_A[6][81] ), .ip2(n9787), .s(n9670), .op(
        n6535) );
  mux2_1 U11310 ( .ip1(\cache_data_A[6][82] ), .ip2(n9788), .s(n9670), .op(
        n6534) );
  mux2_1 U11311 ( .ip1(\cache_data_A[6][83] ), .ip2(n9789), .s(n9670), .op(
        n6533) );
  mux2_1 U11312 ( .ip1(\cache_data_A[6][84] ), .ip2(n9790), .s(n9670), .op(
        n6532) );
  mux2_1 U11313 ( .ip1(\cache_data_A[6][85] ), .ip2(n9791), .s(n9670), .op(
        n6531) );
  mux2_1 U11314 ( .ip1(\cache_data_A[6][86] ), .ip2(n9792), .s(n9670), .op(
        n6530) );
  mux2_1 U11315 ( .ip1(\cache_data_A[6][87] ), .ip2(n9794), .s(n9670), .op(
        n6529) );
  mux2_1 U11316 ( .ip1(\cache_data_A[6][88] ), .ip2(n9795), .s(n9671), .op(
        n6528) );
  mux2_1 U11317 ( .ip1(\cache_data_A[6][89] ), .ip2(n9796), .s(n9671), .op(
        n6527) );
  mux2_1 U11318 ( .ip1(\cache_data_A[6][90] ), .ip2(n9797), .s(n9671), .op(
        n6526) );
  mux2_1 U11319 ( .ip1(\cache_data_A[6][91] ), .ip2(n9798), .s(n9671), .op(
        n6525) );
  mux2_1 U11320 ( .ip1(\cache_data_A[6][92] ), .ip2(n9799), .s(n9671), .op(
        n6524) );
  mux2_1 U11321 ( .ip1(\cache_data_A[6][93] ), .ip2(n9800), .s(n9671), .op(
        n6523) );
  mux2_1 U11322 ( .ip1(\cache_data_A[6][94] ), .ip2(n9801), .s(n9671), .op(
        n6522) );
  mux2_1 U11323 ( .ip1(\cache_data_A[6][95] ), .ip2(n9803), .s(n9671), .op(
        n6521) );
  nor2_1 U11324 ( .ip1(n9762), .ip2(n9672), .op(n9673) );
  mux2_1 U11325 ( .ip1(\cache_data_A[6][96] ), .ip2(n9770), .s(n9673), .op(
        n6520) );
  mux2_1 U11326 ( .ip1(\cache_data_A[6][97] ), .ip2(n9771), .s(n9673), .op(
        n6519) );
  mux2_1 U11327 ( .ip1(\cache_data_A[6][98] ), .ip2(n9772), .s(n9673), .op(
        n6518) );
  mux2_1 U11328 ( .ip1(\cache_data_A[6][99] ), .ip2(n9773), .s(n9673), .op(
        n6517) );
  mux2_1 U11329 ( .ip1(\cache_data_A[6][100] ), .ip2(n9774), .s(n9673), .op(
        n6516) );
  mux2_1 U11330 ( .ip1(\cache_data_A[6][101] ), .ip2(n9775), .s(n9673), .op(
        n6515) );
  mux2_1 U11331 ( .ip1(\cache_data_A[6][102] ), .ip2(n9776), .s(n9673), .op(
        n6514) );
  mux2_1 U11332 ( .ip1(\cache_data_A[6][103] ), .ip2(n9777), .s(n9673), .op(
        n6513) );
  mux2_1 U11333 ( .ip1(\cache_data_A[6][104] ), .ip2(n9778), .s(n9673), .op(
        n6512) );
  buf_1 U11334 ( .ip(n9673), .op(n9674) );
  mux2_1 U11335 ( .ip1(\cache_data_A[6][105] ), .ip2(n9779), .s(n9674), .op(
        n6511) );
  mux2_1 U11336 ( .ip1(\cache_data_A[6][106] ), .ip2(n9780), .s(n9674), .op(
        n6510) );
  mux2_1 U11337 ( .ip1(\cache_data_A[6][107] ), .ip2(n9781), .s(n9673), .op(
        n6509) );
  mux2_1 U11338 ( .ip1(\cache_data_A[6][108] ), .ip2(n9782), .s(n9673), .op(
        n6508) );
  mux2_1 U11339 ( .ip1(\cache_data_A[6][109] ), .ip2(n9783), .s(n9674), .op(
        n6507) );
  mux2_1 U11340 ( .ip1(\cache_data_A[6][110] ), .ip2(n9784), .s(n9673), .op(
        n6506) );
  mux2_1 U11341 ( .ip1(\cache_data_A[6][111] ), .ip2(n9785), .s(n9673), .op(
        n6505) );
  mux2_1 U11342 ( .ip1(\cache_data_A[6][112] ), .ip2(n9786), .s(n9673), .op(
        n6504) );
  mux2_1 U11343 ( .ip1(\cache_data_A[6][113] ), .ip2(n9787), .s(n9673), .op(
        n6503) );
  mux2_1 U11344 ( .ip1(\cache_data_A[6][114] ), .ip2(n9788), .s(n9673), .op(
        n6502) );
  mux2_1 U11345 ( .ip1(\cache_data_A[6][115] ), .ip2(n9789), .s(n9673), .op(
        n6501) );
  mux2_1 U11346 ( .ip1(\cache_data_A[6][116] ), .ip2(n9790), .s(n9673), .op(
        n6500) );
  mux2_1 U11347 ( .ip1(\cache_data_A[6][117] ), .ip2(n9791), .s(n9673), .op(
        n6499) );
  mux2_1 U11348 ( .ip1(\cache_data_A[6][118] ), .ip2(n9792), .s(n9673), .op(
        n6498) );
  mux2_1 U11349 ( .ip1(\cache_data_A[6][119] ), .ip2(n9794), .s(n9673), .op(
        n6497) );
  mux2_1 U11350 ( .ip1(\cache_data_A[6][120] ), .ip2(n9795), .s(n9674), .op(
        n6496) );
  mux2_1 U11351 ( .ip1(\cache_data_A[6][121] ), .ip2(n9796), .s(n9674), .op(
        n6495) );
  mux2_1 U11352 ( .ip1(\cache_data_A[6][122] ), .ip2(n9797), .s(n9674), .op(
        n6494) );
  mux2_1 U11353 ( .ip1(\cache_data_A[6][123] ), .ip2(n9798), .s(n9674), .op(
        n6493) );
  mux2_1 U11354 ( .ip1(\cache_data_A[6][124] ), .ip2(n9799), .s(n9674), .op(
        n6492) );
  mux2_1 U11355 ( .ip1(\cache_data_A[6][125] ), .ip2(n9800), .s(n9674), .op(
        n6491) );
  mux2_1 U11356 ( .ip1(\cache_data_A[6][126] ), .ip2(n9801), .s(n9674), .op(
        n6490) );
  mux2_1 U11357 ( .ip1(\cache_data_A[6][127] ), .ip2(n9803), .s(n9674), .op(
        n6489) );
  nand2_1 U11358 ( .ip1(n9811), .ip2(n9675), .op(n9676) );
  mux2_1 U11359 ( .ip1(n9832), .ip2(\cache_data_A[7][20] ), .s(n9676), .op(
        n6488) );
  mux2_1 U11360 ( .ip1(n9833), .ip2(\cache_data_A[7][21] ), .s(n9676), .op(
        n6487) );
  mux2_1 U11361 ( .ip1(n9835), .ip2(\cache_data_A[7][22] ), .s(n9676), .op(
        n6486) );
  mux2_1 U11362 ( .ip1(n9836), .ip2(\cache_data_A[7][23] ), .s(n9676), .op(
        n6485) );
  mux2_1 U11363 ( .ip1(n9837), .ip2(\cache_data_A[7][24] ), .s(n9676), .op(
        n6484) );
  mux2_1 U11364 ( .ip1(n9838), .ip2(\cache_data_A[7][25] ), .s(n9676), .op(
        n6483) );
  mux2_1 U11365 ( .ip1(n9839), .ip2(\cache_data_A[7][26] ), .s(n9676), .op(
        n6482) );
  mux2_1 U11366 ( .ip1(n9840), .ip2(\cache_data_A[7][27] ), .s(n9676), .op(
        n6481) );
  mux2_1 U11367 ( .ip1(n9841), .ip2(\cache_data_A[7][28] ), .s(n9676), .op(
        n6480) );
  mux2_1 U11368 ( .ip1(n9842), .ip2(\cache_data_A[7][29] ), .s(n9676), .op(
        n6479) );
  mux2_1 U11369 ( .ip1(n9843), .ip2(\cache_data_A[7][30] ), .s(n9676), .op(
        n6478) );
  mux2_1 U11370 ( .ip1(n9845), .ip2(\cache_data_A[7][31] ), .s(n9676), .op(
        n6477) );
  mux2_1 U11371 ( .ip1(n9812), .ip2(\cache_data_A[7][0] ), .s(n9676), .op(
        n6476) );
  mux2_1 U11372 ( .ip1(n9813), .ip2(\cache_data_A[7][1] ), .s(n9676), .op(
        n6475) );
  mux2_1 U11373 ( .ip1(n9814), .ip2(\cache_data_A[7][2] ), .s(n9676), .op(
        n6474) );
  mux2_1 U11374 ( .ip1(n9815), .ip2(\cache_data_A[7][3] ), .s(n9676), .op(
        n6473) );
  mux2_1 U11375 ( .ip1(n9816), .ip2(\cache_data_A[7][4] ), .s(n9676), .op(
        n6472) );
  mux2_1 U11376 ( .ip1(n9817), .ip2(\cache_data_A[7][5] ), .s(n9676), .op(
        n6471) );
  mux2_1 U11377 ( .ip1(n9818), .ip2(\cache_data_A[7][6] ), .s(n9676), .op(
        n6470) );
  buf_1 U11378 ( .ip(n9676), .op(n9677) );
  mux2_1 U11379 ( .ip1(n9819), .ip2(\cache_data_A[7][7] ), .s(n9677), .op(
        n6469) );
  mux2_1 U11380 ( .ip1(n9820), .ip2(\cache_data_A[7][8] ), .s(n9676), .op(
        n6468) );
  mux2_1 U11381 ( .ip1(n9821), .ip2(\cache_data_A[7][9] ), .s(n9677), .op(
        n6467) );
  mux2_1 U11382 ( .ip1(n9822), .ip2(\cache_data_A[7][10] ), .s(n9677), .op(
        n6466) );
  mux2_1 U11383 ( .ip1(n9823), .ip2(\cache_data_A[7][11] ), .s(n9677), .op(
        n6465) );
  mux2_1 U11384 ( .ip1(n9824), .ip2(\cache_data_A[7][12] ), .s(n9677), .op(
        n6464) );
  mux2_1 U11385 ( .ip1(n9825), .ip2(\cache_data_A[7][13] ), .s(n9676), .op(
        n6463) );
  mux2_1 U11386 ( .ip1(n9826), .ip2(\cache_data_A[7][14] ), .s(n9677), .op(
        n6462) );
  mux2_1 U11387 ( .ip1(n9827), .ip2(\cache_data_A[7][15] ), .s(n9677), .op(
        n6461) );
  mux2_1 U11388 ( .ip1(n9828), .ip2(\cache_data_A[7][16] ), .s(n9677), .op(
        n6460) );
  mux2_1 U11389 ( .ip1(n9829), .ip2(\cache_data_A[7][17] ), .s(n9677), .op(
        n6459) );
  mux2_1 U11390 ( .ip1(n9830), .ip2(\cache_data_A[7][18] ), .s(n9677), .op(
        n6458) );
  mux2_1 U11391 ( .ip1(n9831), .ip2(\cache_data_A[7][19] ), .s(n9677), .op(
        n6457) );
  nand2_1 U11392 ( .ip1(n9811), .ip2(n9678), .op(n9679) );
  mux2_1 U11393 ( .ip1(n9770), .ip2(\cache_data_A[7][32] ), .s(n9679), .op(
        n6456) );
  mux2_1 U11394 ( .ip1(n9771), .ip2(\cache_data_A[7][33] ), .s(n9679), .op(
        n6455) );
  mux2_1 U11395 ( .ip1(n9772), .ip2(\cache_data_A[7][34] ), .s(n9679), .op(
        n6454) );
  mux2_1 U11396 ( .ip1(n9773), .ip2(\cache_data_A[7][35] ), .s(n9679), .op(
        n6453) );
  mux2_1 U11397 ( .ip1(n9774), .ip2(\cache_data_A[7][36] ), .s(n9679), .op(
        n6452) );
  mux2_1 U11398 ( .ip1(n9775), .ip2(\cache_data_A[7][37] ), .s(n9679), .op(
        n6451) );
  mux2_1 U11399 ( .ip1(n9776), .ip2(\cache_data_A[7][38] ), .s(n9679), .op(
        n6450) );
  mux2_1 U11400 ( .ip1(n9777), .ip2(\cache_data_A[7][39] ), .s(n9679), .op(
        n6449) );
  mux2_1 U11401 ( .ip1(n9778), .ip2(\cache_data_A[7][40] ), .s(n9679), .op(
        n6448) );
  buf_1 U11402 ( .ip(n9679), .op(n9680) );
  mux2_1 U11403 ( .ip1(n9779), .ip2(\cache_data_A[7][41] ), .s(n9680), .op(
        n6447) );
  mux2_1 U11404 ( .ip1(n9780), .ip2(\cache_data_A[7][42] ), .s(n9679), .op(
        n6446) );
  mux2_1 U11405 ( .ip1(n9781), .ip2(\cache_data_A[7][43] ), .s(n9679), .op(
        n6445) );
  mux2_1 U11406 ( .ip1(n9782), .ip2(\cache_data_A[7][44] ), .s(n9679), .op(
        n6444) );
  mux2_1 U11407 ( .ip1(n9783), .ip2(\cache_data_A[7][45] ), .s(n9679), .op(
        n6443) );
  mux2_1 U11408 ( .ip1(n9784), .ip2(\cache_data_A[7][46] ), .s(n9679), .op(
        n6442) );
  mux2_1 U11409 ( .ip1(n9785), .ip2(\cache_data_A[7][47] ), .s(n9679), .op(
        n6441) );
  mux2_1 U11410 ( .ip1(n9786), .ip2(\cache_data_A[7][48] ), .s(n9679), .op(
        n6440) );
  mux2_1 U11411 ( .ip1(n9787), .ip2(\cache_data_A[7][49] ), .s(n9680), .op(
        n6439) );
  mux2_1 U11412 ( .ip1(n9788), .ip2(\cache_data_A[7][50] ), .s(n9680), .op(
        n6438) );
  mux2_1 U11413 ( .ip1(n9789), .ip2(\cache_data_A[7][51] ), .s(n9680), .op(
        n6437) );
  mux2_1 U11414 ( .ip1(n9832), .ip2(\cache_data_A[7][52] ), .s(n9679), .op(
        n6436) );
  mux2_1 U11415 ( .ip1(n9833), .ip2(\cache_data_A[7][53] ), .s(n9679), .op(
        n6435) );
  mux2_1 U11416 ( .ip1(n9835), .ip2(\cache_data_A[7][54] ), .s(n9679), .op(
        n6434) );
  mux2_1 U11417 ( .ip1(n9836), .ip2(\cache_data_A[7][55] ), .s(n9679), .op(
        n6433) );
  mux2_1 U11418 ( .ip1(n9837), .ip2(\cache_data_A[7][56] ), .s(n9679), .op(
        n6432) );
  mux2_1 U11419 ( .ip1(n9796), .ip2(\cache_data_A[7][57] ), .s(n9680), .op(
        n6431) );
  mux2_1 U11420 ( .ip1(n9797), .ip2(\cache_data_A[7][58] ), .s(n9680), .op(
        n6430) );
  mux2_1 U11421 ( .ip1(n9798), .ip2(\cache_data_A[7][59] ), .s(n9680), .op(
        n6429) );
  mux2_1 U11422 ( .ip1(n9799), .ip2(\cache_data_A[7][60] ), .s(n9680), .op(
        n6428) );
  mux2_1 U11423 ( .ip1(n9800), .ip2(\cache_data_A[7][61] ), .s(n9680), .op(
        n6427) );
  mux2_1 U11424 ( .ip1(n9801), .ip2(\cache_data_A[7][62] ), .s(n9680), .op(
        n6426) );
  mux2_1 U11425 ( .ip1(n9803), .ip2(\cache_data_A[7][63] ), .s(n9680), .op(
        n6425) );
  nor2_1 U11426 ( .ip1(n9769), .ip2(n9681), .op(n9682) );
  mux2_1 U11427 ( .ip1(\cache_data_A[7][64] ), .ip2(n9770), .s(n9682), .op(
        n6424) );
  mux2_1 U11428 ( .ip1(\cache_data_A[7][65] ), .ip2(n9771), .s(n9682), .op(
        n6423) );
  mux2_1 U11429 ( .ip1(\cache_data_A[7][66] ), .ip2(n9772), .s(n9682), .op(
        n6422) );
  mux2_1 U11430 ( .ip1(\cache_data_A[7][67] ), .ip2(n9773), .s(n9682), .op(
        n6421) );
  mux2_1 U11431 ( .ip1(\cache_data_A[7][68] ), .ip2(n9774), .s(n9682), .op(
        n6420) );
  mux2_1 U11432 ( .ip1(\cache_data_A[7][69] ), .ip2(n9775), .s(n9682), .op(
        n6419) );
  mux2_1 U11433 ( .ip1(\cache_data_A[7][70] ), .ip2(n9776), .s(n9682), .op(
        n6418) );
  mux2_1 U11434 ( .ip1(\cache_data_A[7][71] ), .ip2(n9777), .s(n9682), .op(
        n6417) );
  mux2_1 U11435 ( .ip1(\cache_data_A[7][72] ), .ip2(n9778), .s(n9682), .op(
        n6416) );
  buf_1 U11436 ( .ip(n9682), .op(n9683) );
  mux2_1 U11437 ( .ip1(\cache_data_A[7][73] ), .ip2(n9779), .s(n9683), .op(
        n6415) );
  mux2_1 U11438 ( .ip1(\cache_data_A[7][74] ), .ip2(n9780), .s(n9683), .op(
        n6414) );
  mux2_1 U11439 ( .ip1(\cache_data_A[7][75] ), .ip2(n9781), .s(n9682), .op(
        n6413) );
  mux2_1 U11440 ( .ip1(\cache_data_A[7][76] ), .ip2(n9782), .s(n9682), .op(
        n6412) );
  mux2_1 U11441 ( .ip1(\cache_data_A[7][77] ), .ip2(n9783), .s(n9683), .op(
        n6411) );
  mux2_1 U11442 ( .ip1(\cache_data_A[7][78] ), .ip2(n9784), .s(n9682), .op(
        n6410) );
  mux2_1 U11443 ( .ip1(\cache_data_A[7][79] ), .ip2(n9785), .s(n9682), .op(
        n6409) );
  mux2_1 U11444 ( .ip1(\cache_data_A[7][80] ), .ip2(n9786), .s(n9682), .op(
        n6408) );
  mux2_1 U11445 ( .ip1(\cache_data_A[7][81] ), .ip2(n9787), .s(n9682), .op(
        n6407) );
  mux2_1 U11446 ( .ip1(\cache_data_A[7][82] ), .ip2(n9788), .s(n9682), .op(
        n6406) );
  mux2_1 U11447 ( .ip1(\cache_data_A[7][83] ), .ip2(n9789), .s(n9682), .op(
        n6405) );
  mux2_1 U11448 ( .ip1(\cache_data_A[7][84] ), .ip2(n9790), .s(n9682), .op(
        n6404) );
  mux2_1 U11449 ( .ip1(\cache_data_A[7][85] ), .ip2(n9791), .s(n9682), .op(
        n6403) );
  mux2_1 U11450 ( .ip1(\cache_data_A[7][86] ), .ip2(n9792), .s(n9682), .op(
        n6402) );
  mux2_1 U11451 ( .ip1(\cache_data_A[7][87] ), .ip2(n9794), .s(n9682), .op(
        n6401) );
  mux2_1 U11452 ( .ip1(\cache_data_A[7][88] ), .ip2(n9795), .s(n9683), .op(
        n6400) );
  mux2_1 U11453 ( .ip1(\cache_data_A[7][89] ), .ip2(n9796), .s(n9683), .op(
        n6399) );
  mux2_1 U11454 ( .ip1(\cache_data_A[7][90] ), .ip2(n9797), .s(n9683), .op(
        n6398) );
  mux2_1 U11455 ( .ip1(\cache_data_A[7][91] ), .ip2(n9798), .s(n9683), .op(
        n6397) );
  mux2_1 U11456 ( .ip1(\cache_data_A[7][92] ), .ip2(n9799), .s(n9683), .op(
        n6396) );
  mux2_1 U11457 ( .ip1(\cache_data_A[7][93] ), .ip2(n9800), .s(n9683), .op(
        n6395) );
  mux2_1 U11458 ( .ip1(\cache_data_A[7][94] ), .ip2(n9801), .s(n9683), .op(
        n6394) );
  mux2_1 U11459 ( .ip1(\cache_data_A[7][95] ), .ip2(n9803), .s(n9683), .op(
        n6393) );
  nand2_1 U11460 ( .ip1(n9811), .ip2(n9684), .op(n9685) );
  mux2_1 U11461 ( .ip1(n9836), .ip2(\cache_data_A[7][119] ), .s(n9685), .op(
        n6392) );
  mux2_1 U11462 ( .ip1(n9837), .ip2(\cache_data_A[7][120] ), .s(n9685), .op(
        n6391) );
  mux2_1 U11463 ( .ip1(n9796), .ip2(\cache_data_A[7][121] ), .s(n9685), .op(
        n6390) );
  mux2_1 U11464 ( .ip1(n9797), .ip2(\cache_data_A[7][122] ), .s(n9685), .op(
        n6389) );
  mux2_1 U11465 ( .ip1(n9798), .ip2(\cache_data_A[7][123] ), .s(n9685), .op(
        n6388) );
  mux2_1 U11466 ( .ip1(n9799), .ip2(\cache_data_A[7][124] ), .s(n9685), .op(
        n6387) );
  mux2_1 U11467 ( .ip1(n9800), .ip2(\cache_data_A[7][125] ), .s(n9685), .op(
        n6386) );
  mux2_1 U11468 ( .ip1(n9801), .ip2(\cache_data_A[7][126] ), .s(n9685), .op(
        n6385) );
  mux2_1 U11469 ( .ip1(n9803), .ip2(\cache_data_A[7][127] ), .s(n9685), .op(
        n6384) );
  mux2_1 U11470 ( .ip1(n9770), .ip2(\cache_data_A[7][96] ), .s(n9685), .op(
        n6383) );
  mux2_1 U11471 ( .ip1(n9771), .ip2(\cache_data_A[7][97] ), .s(n9685), .op(
        n6382) );
  mux2_1 U11472 ( .ip1(n9772), .ip2(\cache_data_A[7][98] ), .s(n9685), .op(
        n6381) );
  mux2_1 U11473 ( .ip1(n9773), .ip2(\cache_data_A[7][99] ), .s(n9685), .op(
        n6380) );
  mux2_1 U11474 ( .ip1(n9774), .ip2(\cache_data_A[7][100] ), .s(n9685), .op(
        n6379) );
  mux2_1 U11475 ( .ip1(n9775), .ip2(\cache_data_A[7][101] ), .s(n9685), .op(
        n6378) );
  mux2_1 U11476 ( .ip1(n9776), .ip2(\cache_data_A[7][102] ), .s(n9685), .op(
        n6377) );
  buf_1 U11477 ( .ip(n9685), .op(n9686) );
  mux2_1 U11478 ( .ip1(n9777), .ip2(\cache_data_A[7][103] ), .s(n9686), .op(
        n6376) );
  mux2_1 U11479 ( .ip1(n9778), .ip2(\cache_data_A[7][104] ), .s(n9685), .op(
        n6375) );
  mux2_1 U11480 ( .ip1(n9779), .ip2(\cache_data_A[7][105] ), .s(n9685), .op(
        n6374) );
  mux2_1 U11481 ( .ip1(n9780), .ip2(\cache_data_A[7][106] ), .s(n9685), .op(
        n6373) );
  mux2_1 U11482 ( .ip1(n9781), .ip2(\cache_data_A[7][107] ), .s(n9686), .op(
        n6372) );
  mux2_1 U11483 ( .ip1(n9782), .ip2(\cache_data_A[7][108] ), .s(n9685), .op(
        n6371) );
  mux2_1 U11484 ( .ip1(n9783), .ip2(\cache_data_A[7][109] ), .s(n9686), .op(
        n6370) );
  mux2_1 U11485 ( .ip1(n9784), .ip2(\cache_data_A[7][110] ), .s(n9686), .op(
        n6369) );
  mux2_1 U11486 ( .ip1(n9785), .ip2(\cache_data_A[7][111] ), .s(n9685), .op(
        n6368) );
  mux2_1 U11487 ( .ip1(n9786), .ip2(\cache_data_A[7][112] ), .s(n9686), .op(
        n6367) );
  mux2_1 U11488 ( .ip1(n9787), .ip2(\cache_data_A[7][113] ), .s(n9686), .op(
        n6366) );
  mux2_1 U11489 ( .ip1(n9788), .ip2(\cache_data_A[7][114] ), .s(n9686), .op(
        n6365) );
  mux2_1 U11490 ( .ip1(n9789), .ip2(\cache_data_A[7][115] ), .s(n9686), .op(
        n6364) );
  mux2_1 U11491 ( .ip1(n9790), .ip2(\cache_data_A[7][116] ), .s(n9686), .op(
        n6363) );
  mux2_1 U11492 ( .ip1(n9833), .ip2(\cache_data_A[7][117] ), .s(n9686), .op(
        n6362) );
  mux2_1 U11493 ( .ip1(n9835), .ip2(\cache_data_A[7][118] ), .s(n9686), .op(
        n6361) );
  nand3_1 U11494 ( .ip1(n9885), .ip2(n9687), .ip3(n9846), .op(n9689) );
  nor3_1 U11495 ( .ip1(mem_data_cnt[3]), .ip2(mem_data_cnt[2]), .ip3(n9702), 
        .op(n13170) );
  nand2_1 U11496 ( .ip1(n9703), .ip2(n13170), .op(n9688) );
  nand2_1 U11497 ( .ip1(n9689), .ip2(n9688), .op(n9756) );
  nand2_1 U11498 ( .ip1(n13293), .ip2(n9756), .op(n9768) );
  nor2_1 U11499 ( .ip1(n9860), .ip2(n9768), .op(n9690) );
  buf_1 U11500 ( .ip(n9690), .op(n9691) );
  mux2_1 U11501 ( .ip1(\cache_data_B[0][0] ), .ip2(n9770), .s(n9691), .op(
        n6360) );
  mux2_1 U11502 ( .ip1(\cache_data_B[0][1] ), .ip2(n9771), .s(n9690), .op(
        n6359) );
  mux2_1 U11503 ( .ip1(\cache_data_B[0][2] ), .ip2(n9772), .s(n9690), .op(
        n6358) );
  mux2_1 U11504 ( .ip1(\cache_data_B[0][3] ), .ip2(n9773), .s(n9690), .op(
        n6357) );
  mux2_1 U11505 ( .ip1(\cache_data_B[0][4] ), .ip2(n9774), .s(n9690), .op(
        n6356) );
  mux2_1 U11506 ( .ip1(\cache_data_B[0][5] ), .ip2(n9775), .s(n9690), .op(
        n6355) );
  mux2_1 U11507 ( .ip1(\cache_data_B[0][6] ), .ip2(n9776), .s(n9690), .op(
        n6354) );
  mux2_1 U11508 ( .ip1(\cache_data_B[0][7] ), .ip2(n9777), .s(n9690), .op(
        n6353) );
  mux2_1 U11509 ( .ip1(\cache_data_B[0][8] ), .ip2(n9778), .s(n9690), .op(
        n6352) );
  mux2_1 U11510 ( .ip1(\cache_data_B[0][9] ), .ip2(n9779), .s(n9691), .op(
        n6351) );
  mux2_1 U11511 ( .ip1(\cache_data_B[0][10] ), .ip2(n9780), .s(n9691), .op(
        n6350) );
  mux2_1 U11512 ( .ip1(\cache_data_B[0][11] ), .ip2(n9781), .s(n9690), .op(
        n6349) );
  mux2_1 U11513 ( .ip1(\cache_data_B[0][12] ), .ip2(n9782), .s(n9690), .op(
        n6348) );
  mux2_1 U11514 ( .ip1(\cache_data_B[0][13] ), .ip2(n9783), .s(n9690), .op(
        n6347) );
  mux2_1 U11515 ( .ip1(\cache_data_B[0][14] ), .ip2(n9784), .s(n9690), .op(
        n6346) );
  mux2_1 U11516 ( .ip1(\cache_data_B[0][15] ), .ip2(n9785), .s(n9690), .op(
        n6345) );
  mux2_1 U11517 ( .ip1(\cache_data_B[0][16] ), .ip2(n9786), .s(n9690), .op(
        n6344) );
  mux2_1 U11518 ( .ip1(\cache_data_B[0][17] ), .ip2(n9787), .s(n9690), .op(
        n6343) );
  mux2_1 U11519 ( .ip1(\cache_data_B[0][18] ), .ip2(n9788), .s(n9690), .op(
        n6342) );
  mux2_1 U11520 ( .ip1(\cache_data_B[0][19] ), .ip2(n9789), .s(n9690), .op(
        n6341) );
  mux2_1 U11521 ( .ip1(\cache_data_B[0][20] ), .ip2(n9790), .s(n9690), .op(
        n6340) );
  mux2_1 U11522 ( .ip1(\cache_data_B[0][21] ), .ip2(n9791), .s(n9690), .op(
        n6339) );
  mux2_1 U11523 ( .ip1(\cache_data_B[0][22] ), .ip2(n9792), .s(n9690), .op(
        n6338) );
  mux2_1 U11524 ( .ip1(\cache_data_B[0][23] ), .ip2(n9794), .s(n9690), .op(
        n6337) );
  mux2_1 U11525 ( .ip1(\cache_data_B[0][24] ), .ip2(n9795), .s(n9691), .op(
        n6336) );
  mux2_1 U11526 ( .ip1(\cache_data_B[0][25] ), .ip2(n9796), .s(n9691), .op(
        n6335) );
  mux2_1 U11527 ( .ip1(\cache_data_B[0][26] ), .ip2(n9797), .s(n9691), .op(
        n6334) );
  mux2_1 U11528 ( .ip1(\cache_data_B[0][27] ), .ip2(n9798), .s(n9691), .op(
        n6333) );
  mux2_1 U11529 ( .ip1(\cache_data_B[0][28] ), .ip2(n9799), .s(n9691), .op(
        n6332) );
  mux2_1 U11530 ( .ip1(\cache_data_B[0][29] ), .ip2(n9800), .s(n9691), .op(
        n6331) );
  mux2_1 U11531 ( .ip1(\cache_data_B[0][30] ), .ip2(n9801), .s(n9691), .op(
        n6330) );
  mux2_1 U11532 ( .ip1(\cache_data_B[0][31] ), .ip2(n9803), .s(n9691), .op(
        n6329) );
  nor3_1 U11533 ( .ip1(mem_data_cnt[3]), .ip2(n9702), .ip3(n9700), .op(n13182)
         );
  nand2_1 U11534 ( .ip1(n13182), .ip2(n9703), .op(n9693) );
  nor3_1 U11535 ( .ip1(addr_resp[3]), .ip2(n9925), .ip3(n9705), .op(n12563) );
  nand2_1 U11536 ( .ip1(n12563), .ip2(n9846), .op(n9692) );
  nand2_1 U11537 ( .ip1(n9693), .ip2(n9692), .op(n9804) );
  nand2_1 U11538 ( .ip1(n9708), .ip2(n9804), .op(n9694) );
  mux2_1 U11539 ( .ip1(n9770), .ip2(\cache_data_B[0][32] ), .s(n9694), .op(
        n6328) );
  mux2_1 U11540 ( .ip1(n9771), .ip2(\cache_data_B[0][33] ), .s(n9694), .op(
        n6327) );
  mux2_1 U11541 ( .ip1(n9772), .ip2(\cache_data_B[0][34] ), .s(n9694), .op(
        n6326) );
  mux2_1 U11542 ( .ip1(n9773), .ip2(\cache_data_B[0][35] ), .s(n9694), .op(
        n6325) );
  mux2_1 U11543 ( .ip1(n9774), .ip2(\cache_data_B[0][36] ), .s(n9694), .op(
        n6324) );
  mux2_1 U11544 ( .ip1(n9775), .ip2(\cache_data_B[0][37] ), .s(n9694), .op(
        n6323) );
  mux2_1 U11545 ( .ip1(n9776), .ip2(\cache_data_B[0][38] ), .s(n9694), .op(
        n6322) );
  mux2_1 U11546 ( .ip1(n9777), .ip2(\cache_data_B[0][39] ), .s(n9694), .op(
        n6321) );
  mux2_1 U11547 ( .ip1(n9778), .ip2(\cache_data_B[0][40] ), .s(n9694), .op(
        n6320) );
  mux2_1 U11548 ( .ip1(n9779), .ip2(\cache_data_B[0][41] ), .s(n9694), .op(
        n6319) );
  mux2_1 U11549 ( .ip1(n9780), .ip2(\cache_data_B[0][42] ), .s(n9694), .op(
        n6318) );
  buf_1 U11550 ( .ip(n9694), .op(n9695) );
  mux2_1 U11551 ( .ip1(n9781), .ip2(\cache_data_B[0][43] ), .s(n9695), .op(
        n6317) );
  mux2_1 U11552 ( .ip1(n9782), .ip2(\cache_data_B[0][44] ), .s(n9694), .op(
        n6316) );
  mux2_1 U11553 ( .ip1(n9783), .ip2(\cache_data_B[0][45] ), .s(n9694), .op(
        n6315) );
  mux2_1 U11554 ( .ip1(n9784), .ip2(\cache_data_B[0][46] ), .s(n9694), .op(
        n6314) );
  mux2_1 U11555 ( .ip1(n9785), .ip2(\cache_data_B[0][47] ), .s(n9694), .op(
        n6313) );
  mux2_1 U11556 ( .ip1(n9786), .ip2(\cache_data_B[0][48] ), .s(n9695), .op(
        n6312) );
  mux2_1 U11557 ( .ip1(n9787), .ip2(\cache_data_B[0][49] ), .s(n9694), .op(
        n6311) );
  mux2_1 U11558 ( .ip1(n9788), .ip2(\cache_data_B[0][50] ), .s(n9694), .op(
        n6310) );
  mux2_1 U11559 ( .ip1(n9789), .ip2(\cache_data_B[0][51] ), .s(n9694), .op(
        n6309) );
  mux2_1 U11560 ( .ip1(n9832), .ip2(\cache_data_B[0][52] ), .s(n9694), .op(
        n6308) );
  mux2_1 U11561 ( .ip1(n9791), .ip2(\cache_data_B[0][53] ), .s(n9695), .op(
        n6307) );
  mux2_1 U11562 ( .ip1(n9792), .ip2(\cache_data_B[0][54] ), .s(n9694), .op(
        n6306) );
  mux2_1 U11563 ( .ip1(n9794), .ip2(\cache_data_B[0][55] ), .s(n9694), .op(
        n6305) );
  mux2_1 U11564 ( .ip1(n9795), .ip2(\cache_data_B[0][56] ), .s(n9695), .op(
        n6304) );
  mux2_1 U11565 ( .ip1(n9796), .ip2(\cache_data_B[0][57] ), .s(n9695), .op(
        n6303) );
  mux2_1 U11566 ( .ip1(n9797), .ip2(\cache_data_B[0][58] ), .s(n9695), .op(
        n6302) );
  mux2_1 U11567 ( .ip1(n9798), .ip2(\cache_data_B[0][59] ), .s(n9695), .op(
        n6301) );
  mux2_1 U11568 ( .ip1(n9799), .ip2(\cache_data_B[0][60] ), .s(n9695), .op(
        n6300) );
  mux2_1 U11569 ( .ip1(n9800), .ip2(\cache_data_B[0][61] ), .s(n9695), .op(
        n6299) );
  mux2_1 U11570 ( .ip1(n9801), .ip2(\cache_data_B[0][62] ), .s(n9695), .op(
        n6298) );
  mux2_1 U11571 ( .ip1(n9803), .ip2(\cache_data_B[0][63] ), .s(n9695), .op(
        n6297) );
  nand3_1 U11572 ( .ip1(n9885), .ip2(n9846), .ip3(n9905), .op(n9697) );
  nor3_1 U11573 ( .ip1(mem_data_cnt[2]), .ip2(n9701), .ip3(n9702), .op(n13168)
         );
  nand2_1 U11574 ( .ip1(n9703), .ip2(n13168), .op(n9696) );
  nand2_1 U11575 ( .ip1(n9697), .ip2(n9696), .op(n9807) );
  nand2_1 U11576 ( .ip1(n9708), .ip2(n9807), .op(n9698) );
  mux2_1 U11577 ( .ip1(n9795), .ip2(\cache_data_B[0][88] ), .s(n9698), .op(
        n6296) );
  mux2_1 U11578 ( .ip1(n9796), .ip2(\cache_data_B[0][89] ), .s(n9698), .op(
        n6295) );
  mux2_1 U11579 ( .ip1(n9797), .ip2(\cache_data_B[0][90] ), .s(n9698), .op(
        n6294) );
  mux2_1 U11580 ( .ip1(n9798), .ip2(\cache_data_B[0][91] ), .s(n9698), .op(
        n6293) );
  mux2_1 U11581 ( .ip1(n9799), .ip2(\cache_data_B[0][92] ), .s(n9698), .op(
        n6292) );
  mux2_1 U11582 ( .ip1(n9800), .ip2(\cache_data_B[0][93] ), .s(n9698), .op(
        n6291) );
  mux2_1 U11583 ( .ip1(n9801), .ip2(\cache_data_B[0][94] ), .s(n9698), .op(
        n6290) );
  mux2_1 U11584 ( .ip1(n9803), .ip2(\cache_data_B[0][95] ), .s(n9698), .op(
        n6289) );
  mux2_1 U11585 ( .ip1(n9770), .ip2(\cache_data_B[0][64] ), .s(n9698), .op(
        n6288) );
  mux2_1 U11586 ( .ip1(n9771), .ip2(\cache_data_B[0][65] ), .s(n9698), .op(
        n6287) );
  buf_1 U11587 ( .ip(n9698), .op(n9699) );
  mux2_1 U11588 ( .ip1(n9772), .ip2(\cache_data_B[0][66] ), .s(n9699), .op(
        n6286) );
  mux2_1 U11589 ( .ip1(n9773), .ip2(\cache_data_B[0][67] ), .s(n9698), .op(
        n6285) );
  mux2_1 U11590 ( .ip1(n9774), .ip2(\cache_data_B[0][68] ), .s(n9698), .op(
        n6284) );
  mux2_1 U11591 ( .ip1(n9775), .ip2(\cache_data_B[0][69] ), .s(n9698), .op(
        n6283) );
  mux2_1 U11592 ( .ip1(n9776), .ip2(\cache_data_B[0][70] ), .s(n9698), .op(
        n6282) );
  mux2_1 U11593 ( .ip1(n9777), .ip2(\cache_data_B[0][71] ), .s(n9698), .op(
        n6281) );
  mux2_1 U11594 ( .ip1(n9778), .ip2(\cache_data_B[0][72] ), .s(n9698), .op(
        n6280) );
  mux2_1 U11595 ( .ip1(n9779), .ip2(\cache_data_B[0][73] ), .s(n9698), .op(
        n6279) );
  mux2_1 U11596 ( .ip1(n9780), .ip2(\cache_data_B[0][74] ), .s(n9698), .op(
        n6278) );
  mux2_1 U11597 ( .ip1(n9781), .ip2(\cache_data_B[0][75] ), .s(n9698), .op(
        n6277) );
  mux2_1 U11598 ( .ip1(n9782), .ip2(\cache_data_B[0][76] ), .s(n9698), .op(
        n6276) );
  mux2_1 U11599 ( .ip1(n9783), .ip2(\cache_data_B[0][77] ), .s(n9698), .op(
        n6275) );
  mux2_1 U11600 ( .ip1(n9784), .ip2(\cache_data_B[0][78] ), .s(n9699), .op(
        n6274) );
  mux2_1 U11601 ( .ip1(n9785), .ip2(\cache_data_B[0][79] ), .s(n9699), .op(
        n6273) );
  mux2_1 U11602 ( .ip1(n9786), .ip2(\cache_data_B[0][80] ), .s(n9699), .op(
        n6272) );
  mux2_1 U11603 ( .ip1(n9787), .ip2(\cache_data_B[0][81] ), .s(n9699), .op(
        n6271) );
  mux2_1 U11604 ( .ip1(n9788), .ip2(\cache_data_B[0][82] ), .s(n9699), .op(
        n6270) );
  mux2_1 U11605 ( .ip1(n9831), .ip2(\cache_data_B[0][83] ), .s(n9699), .op(
        n6269) );
  mux2_1 U11606 ( .ip1(n9790), .ip2(\cache_data_B[0][84] ), .s(n9699), .op(
        n6268) );
  mux2_1 U11607 ( .ip1(n9791), .ip2(\cache_data_B[0][85] ), .s(n9699), .op(
        n6267) );
  mux2_1 U11608 ( .ip1(n9835), .ip2(\cache_data_B[0][86] ), .s(n9699), .op(
        n6266) );
  mux2_1 U11609 ( .ip1(n9836), .ip2(\cache_data_B[0][87] ), .s(n9699), .op(
        n6265) );
  nor3_1 U11610 ( .ip1(n9702), .ip2(n9701), .ip3(n9700), .op(n13166) );
  nand2_1 U11611 ( .ip1(n13166), .ip2(n9703), .op(n9707) );
  nor3_1 U11612 ( .ip1(n9925), .ip2(n9705), .ip3(n9704), .op(n12573) );
  nand2_1 U11613 ( .ip1(n12573), .ip2(n9846), .op(n9706) );
  nand2_1 U11614 ( .ip1(n9707), .ip2(n9706), .op(n9810) );
  nand2_1 U11615 ( .ip1(n9708), .ip2(n9810), .op(n9709) );
  mux2_1 U11616 ( .ip1(n9770), .ip2(\cache_data_B[0][96] ), .s(n9709), .op(
        n6264) );
  buf_1 U11617 ( .ip(n9709), .op(n9710) );
  mux2_1 U11618 ( .ip1(n9771), .ip2(\cache_data_B[0][97] ), .s(n9710), .op(
        n6263) );
  mux2_1 U11619 ( .ip1(n9772), .ip2(\cache_data_B[0][98] ), .s(n9709), .op(
        n6262) );
  mux2_1 U11620 ( .ip1(n9773), .ip2(\cache_data_B[0][99] ), .s(n9709), .op(
        n6261) );
  mux2_1 U11621 ( .ip1(n9774), .ip2(\cache_data_B[0][100] ), .s(n9709), .op(
        n6260) );
  mux2_1 U11622 ( .ip1(n9775), .ip2(\cache_data_B[0][101] ), .s(n9709), .op(
        n6259) );
  mux2_1 U11623 ( .ip1(n9776), .ip2(\cache_data_B[0][102] ), .s(n9709), .op(
        n6258) );
  mux2_1 U11624 ( .ip1(n9777), .ip2(\cache_data_B[0][103] ), .s(n9709), .op(
        n6257) );
  mux2_1 U11625 ( .ip1(n9778), .ip2(\cache_data_B[0][104] ), .s(n9709), .op(
        n6256) );
  mux2_1 U11626 ( .ip1(n9779), .ip2(\cache_data_B[0][105] ), .s(n9709), .op(
        n6255) );
  mux2_1 U11627 ( .ip1(n9780), .ip2(\cache_data_B[0][106] ), .s(n9709), .op(
        n6254) );
  mux2_1 U11628 ( .ip1(n9781), .ip2(\cache_data_B[0][107] ), .s(n9709), .op(
        n6253) );
  mux2_1 U11629 ( .ip1(n9782), .ip2(\cache_data_B[0][108] ), .s(n9709), .op(
        n6252) );
  mux2_1 U11630 ( .ip1(n9783), .ip2(\cache_data_B[0][109] ), .s(n9709), .op(
        n6251) );
  mux2_1 U11631 ( .ip1(n9784), .ip2(\cache_data_B[0][110] ), .s(n9710), .op(
        n6250) );
  mux2_1 U11632 ( .ip1(n9785), .ip2(\cache_data_B[0][111] ), .s(n9709), .op(
        n6249) );
  mux2_1 U11633 ( .ip1(n9786), .ip2(\cache_data_B[0][112] ), .s(n9710), .op(
        n6248) );
  mux2_1 U11634 ( .ip1(n9787), .ip2(\cache_data_B[0][113] ), .s(n9710), .op(
        n6247) );
  mux2_1 U11635 ( .ip1(n9788), .ip2(\cache_data_B[0][114] ), .s(n9709), .op(
        n6246) );
  mux2_1 U11636 ( .ip1(n9789), .ip2(\cache_data_B[0][115] ), .s(n9709), .op(
        n6245) );
  mux2_1 U11637 ( .ip1(n9832), .ip2(\cache_data_B[0][116] ), .s(n9709), .op(
        n6244) );
  mux2_1 U11638 ( .ip1(n9833), .ip2(\cache_data_B[0][117] ), .s(n9709), .op(
        n6243) );
  mux2_1 U11639 ( .ip1(n9792), .ip2(\cache_data_B[0][118] ), .s(n9709), .op(
        n6242) );
  mux2_1 U11640 ( .ip1(n9836), .ip2(\cache_data_B[0][119] ), .s(n9710), .op(
        n6241) );
  mux2_1 U11641 ( .ip1(n9837), .ip2(\cache_data_B[0][120] ), .s(n9709), .op(
        n6240) );
  mux2_1 U11642 ( .ip1(n9796), .ip2(\cache_data_B[0][121] ), .s(n9709), .op(
        n6239) );
  mux2_1 U11643 ( .ip1(n9797), .ip2(\cache_data_B[0][122] ), .s(n9710), .op(
        n6238) );
  mux2_1 U11644 ( .ip1(n9798), .ip2(\cache_data_B[0][123] ), .s(n9710), .op(
        n6237) );
  mux2_1 U11645 ( .ip1(n9799), .ip2(\cache_data_B[0][124] ), .s(n9710), .op(
        n6236) );
  mux2_1 U11646 ( .ip1(n9800), .ip2(\cache_data_B[0][125] ), .s(n9710), .op(
        n6235) );
  mux2_1 U11647 ( .ip1(n9801), .ip2(\cache_data_B[0][126] ), .s(n9710), .op(
        n6234) );
  mux2_1 U11648 ( .ip1(n9803), .ip2(\cache_data_B[0][127] ), .s(n9710), .op(
        n6233) );
  nor2_1 U11649 ( .ip1(n9862), .ip2(n9768), .op(n9711) );
  buf_1 U11650 ( .ip(n9711), .op(n9712) );
  mux2_1 U11651 ( .ip1(\cache_data_B[1][0] ), .ip2(n9770), .s(n9712), .op(
        n6232) );
  mux2_1 U11652 ( .ip1(\cache_data_B[1][1] ), .ip2(n9771), .s(n9711), .op(
        n6231) );
  mux2_1 U11653 ( .ip1(\cache_data_B[1][2] ), .ip2(n9772), .s(n9711), .op(
        n6230) );
  mux2_1 U11654 ( .ip1(\cache_data_B[1][3] ), .ip2(n9773), .s(n9711), .op(
        n6229) );
  mux2_1 U11655 ( .ip1(\cache_data_B[1][4] ), .ip2(n9774), .s(n9711), .op(
        n6228) );
  mux2_1 U11656 ( .ip1(\cache_data_B[1][5] ), .ip2(n9775), .s(n9711), .op(
        n6227) );
  mux2_1 U11657 ( .ip1(\cache_data_B[1][6] ), .ip2(n9776), .s(n9711), .op(
        n6226) );
  mux2_1 U11658 ( .ip1(\cache_data_B[1][7] ), .ip2(n9777), .s(n9711), .op(
        n6225) );
  mux2_1 U11659 ( .ip1(\cache_data_B[1][8] ), .ip2(n9778), .s(n9711), .op(
        n6224) );
  mux2_1 U11660 ( .ip1(\cache_data_B[1][9] ), .ip2(n9779), .s(n9712), .op(
        n6223) );
  mux2_1 U11661 ( .ip1(\cache_data_B[1][10] ), .ip2(n9780), .s(n9712), .op(
        n6222) );
  mux2_1 U11662 ( .ip1(\cache_data_B[1][11] ), .ip2(n9781), .s(n9711), .op(
        n6221) );
  mux2_1 U11663 ( .ip1(\cache_data_B[1][12] ), .ip2(n9782), .s(n9711), .op(
        n6220) );
  mux2_1 U11664 ( .ip1(\cache_data_B[1][13] ), .ip2(n9783), .s(n9711), .op(
        n6219) );
  mux2_1 U11665 ( .ip1(\cache_data_B[1][14] ), .ip2(n9784), .s(n9711), .op(
        n6218) );
  mux2_1 U11666 ( .ip1(\cache_data_B[1][15] ), .ip2(n9785), .s(n9711), .op(
        n6217) );
  mux2_1 U11667 ( .ip1(\cache_data_B[1][16] ), .ip2(n9786), .s(n9711), .op(
        n6216) );
  mux2_1 U11668 ( .ip1(\cache_data_B[1][17] ), .ip2(n9787), .s(n9711), .op(
        n6215) );
  mux2_1 U11669 ( .ip1(\cache_data_B[1][18] ), .ip2(n9788), .s(n9711), .op(
        n6214) );
  mux2_1 U11670 ( .ip1(\cache_data_B[1][19] ), .ip2(n9789), .s(n9711), .op(
        n6213) );
  mux2_1 U11671 ( .ip1(\cache_data_B[1][20] ), .ip2(n9790), .s(n9711), .op(
        n6212) );
  mux2_1 U11672 ( .ip1(\cache_data_B[1][21] ), .ip2(n9791), .s(n9711), .op(
        n6211) );
  mux2_1 U11673 ( .ip1(\cache_data_B[1][22] ), .ip2(n9792), .s(n9711), .op(
        n6210) );
  mux2_1 U11674 ( .ip1(\cache_data_B[1][23] ), .ip2(n9794), .s(n9711), .op(
        n6209) );
  mux2_1 U11675 ( .ip1(\cache_data_B[1][24] ), .ip2(n9795), .s(n9712), .op(
        n6208) );
  mux2_1 U11676 ( .ip1(\cache_data_B[1][25] ), .ip2(n9796), .s(n9712), .op(
        n6207) );
  mux2_1 U11677 ( .ip1(\cache_data_B[1][26] ), .ip2(n9797), .s(n9712), .op(
        n6206) );
  mux2_1 U11678 ( .ip1(\cache_data_B[1][27] ), .ip2(n9798), .s(n9712), .op(
        n6205) );
  mux2_1 U11679 ( .ip1(\cache_data_B[1][28] ), .ip2(n9799), .s(n9712), .op(
        n6204) );
  mux2_1 U11680 ( .ip1(\cache_data_B[1][29] ), .ip2(n9800), .s(n9712), .op(
        n6203) );
  mux2_1 U11681 ( .ip1(\cache_data_B[1][30] ), .ip2(n9801), .s(n9712), .op(
        n6202) );
  mux2_1 U11682 ( .ip1(\cache_data_B[1][31] ), .ip2(n9803), .s(n9712), .op(
        n6201) );
  nand2_1 U11683 ( .ip1(n9717), .ip2(n9804), .op(n9713) );
  mux2_1 U11684 ( .ip1(n9798), .ip2(\cache_data_B[1][59] ), .s(n9713), .op(
        n6200) );
  mux2_1 U11685 ( .ip1(n9799), .ip2(\cache_data_B[1][60] ), .s(n9713), .op(
        n6199) );
  mux2_1 U11686 ( .ip1(n9800), .ip2(\cache_data_B[1][61] ), .s(n9713), .op(
        n6198) );
  mux2_1 U11687 ( .ip1(n9801), .ip2(\cache_data_B[1][62] ), .s(n9713), .op(
        n6197) );
  mux2_1 U11688 ( .ip1(n9803), .ip2(\cache_data_B[1][63] ), .s(n9713), .op(
        n6196) );
  mux2_1 U11689 ( .ip1(n9770), .ip2(\cache_data_B[1][32] ), .s(n9713), .op(
        n6195) );
  mux2_1 U11690 ( .ip1(n9771), .ip2(\cache_data_B[1][33] ), .s(n9713), .op(
        n6194) );
  mux2_1 U11691 ( .ip1(n9772), .ip2(\cache_data_B[1][34] ), .s(n9713), .op(
        n6193) );
  mux2_1 U11692 ( .ip1(n9773), .ip2(\cache_data_B[1][35] ), .s(n9713), .op(
        n6192) );
  buf_1 U11693 ( .ip(n9713), .op(n9714) );
  mux2_1 U11694 ( .ip1(n9774), .ip2(\cache_data_B[1][36] ), .s(n9714), .op(
        n6191) );
  mux2_1 U11695 ( .ip1(n9775), .ip2(\cache_data_B[1][37] ), .s(n9713), .op(
        n6190) );
  mux2_1 U11696 ( .ip1(n9776), .ip2(\cache_data_B[1][38] ), .s(n9713), .op(
        n6189) );
  mux2_1 U11697 ( .ip1(n9777), .ip2(\cache_data_B[1][39] ), .s(n9713), .op(
        n6188) );
  mux2_1 U11698 ( .ip1(n9778), .ip2(\cache_data_B[1][40] ), .s(n9713), .op(
        n6187) );
  mux2_1 U11699 ( .ip1(n9779), .ip2(\cache_data_B[1][41] ), .s(n9713), .op(
        n6186) );
  mux2_1 U11700 ( .ip1(n9780), .ip2(\cache_data_B[1][42] ), .s(n9713), .op(
        n6185) );
  mux2_1 U11701 ( .ip1(n9781), .ip2(\cache_data_B[1][43] ), .s(n9713), .op(
        n6184) );
  mux2_1 U11702 ( .ip1(n9782), .ip2(\cache_data_B[1][44] ), .s(n9713), .op(
        n6183) );
  mux2_1 U11703 ( .ip1(n9783), .ip2(\cache_data_B[1][45] ), .s(n9713), .op(
        n6182) );
  mux2_1 U11704 ( .ip1(n9784), .ip2(\cache_data_B[1][46] ), .s(n9713), .op(
        n6181) );
  mux2_1 U11705 ( .ip1(n9785), .ip2(\cache_data_B[1][47] ), .s(n9714), .op(
        n6180) );
  mux2_1 U11706 ( .ip1(n9786), .ip2(\cache_data_B[1][48] ), .s(n9713), .op(
        n6179) );
  mux2_1 U11707 ( .ip1(n9787), .ip2(\cache_data_B[1][49] ), .s(n9713), .op(
        n6178) );
  mux2_1 U11708 ( .ip1(n9788), .ip2(\cache_data_B[1][50] ), .s(n9714), .op(
        n6177) );
  mux2_1 U11709 ( .ip1(n9831), .ip2(\cache_data_B[1][51] ), .s(n9714), .op(
        n6176) );
  mux2_1 U11710 ( .ip1(n9790), .ip2(\cache_data_B[1][52] ), .s(n9714), .op(
        n6175) );
  mux2_1 U11711 ( .ip1(n9791), .ip2(\cache_data_B[1][53] ), .s(n9714), .op(
        n6174) );
  mux2_1 U11712 ( .ip1(n9792), .ip2(\cache_data_B[1][54] ), .s(n9714), .op(
        n6173) );
  mux2_1 U11713 ( .ip1(n9794), .ip2(\cache_data_B[1][55] ), .s(n9714), .op(
        n6172) );
  mux2_1 U11714 ( .ip1(n9795), .ip2(\cache_data_B[1][56] ), .s(n9714), .op(
        n6171) );
  mux2_1 U11715 ( .ip1(n9796), .ip2(\cache_data_B[1][57] ), .s(n9714), .op(
        n6170) );
  mux2_1 U11716 ( .ip1(n9797), .ip2(\cache_data_B[1][58] ), .s(n9714), .op(
        n6169) );
  nand2_1 U11717 ( .ip1(n13293), .ip2(n9807), .op(n9761) );
  nor2_1 U11718 ( .ip1(n9862), .ip2(n9761), .op(n9715) );
  buf_1 U11719 ( .ip(n9715), .op(n9716) );
  mux2_1 U11720 ( .ip1(\cache_data_B[1][64] ), .ip2(n9770), .s(n9716), .op(
        n6168) );
  mux2_1 U11721 ( .ip1(\cache_data_B[1][65] ), .ip2(n9771), .s(n9715), .op(
        n6167) );
  mux2_1 U11722 ( .ip1(\cache_data_B[1][66] ), .ip2(n9772), .s(n9715), .op(
        n6166) );
  mux2_1 U11723 ( .ip1(\cache_data_B[1][67] ), .ip2(n9773), .s(n9715), .op(
        n6165) );
  mux2_1 U11724 ( .ip1(\cache_data_B[1][68] ), .ip2(n9774), .s(n9715), .op(
        n6164) );
  mux2_1 U11725 ( .ip1(\cache_data_B[1][69] ), .ip2(n9775), .s(n9715), .op(
        n6163) );
  mux2_1 U11726 ( .ip1(\cache_data_B[1][70] ), .ip2(n9776), .s(n9715), .op(
        n6162) );
  mux2_1 U11727 ( .ip1(\cache_data_B[1][71] ), .ip2(n9777), .s(n9715), .op(
        n6161) );
  mux2_1 U11728 ( .ip1(\cache_data_B[1][72] ), .ip2(n9778), .s(n9715), .op(
        n6160) );
  mux2_1 U11729 ( .ip1(\cache_data_B[1][73] ), .ip2(n9779), .s(n9716), .op(
        n6159) );
  mux2_1 U11730 ( .ip1(\cache_data_B[1][74] ), .ip2(n9780), .s(n9716), .op(
        n6158) );
  mux2_1 U11731 ( .ip1(\cache_data_B[1][75] ), .ip2(n9781), .s(n9715), .op(
        n6157) );
  mux2_1 U11732 ( .ip1(\cache_data_B[1][76] ), .ip2(n9782), .s(n9715), .op(
        n6156) );
  mux2_1 U11733 ( .ip1(\cache_data_B[1][77] ), .ip2(n9783), .s(n9715), .op(
        n6155) );
  mux2_1 U11734 ( .ip1(\cache_data_B[1][78] ), .ip2(n9784), .s(n9715), .op(
        n6154) );
  mux2_1 U11735 ( .ip1(\cache_data_B[1][79] ), .ip2(n9785), .s(n9715), .op(
        n6153) );
  mux2_1 U11736 ( .ip1(\cache_data_B[1][80] ), .ip2(n9786), .s(n9715), .op(
        n6152) );
  mux2_1 U11737 ( .ip1(\cache_data_B[1][81] ), .ip2(n9787), .s(n9715), .op(
        n6151) );
  mux2_1 U11738 ( .ip1(\cache_data_B[1][82] ), .ip2(n9788), .s(n9715), .op(
        n6150) );
  mux2_1 U11739 ( .ip1(\cache_data_B[1][83] ), .ip2(n9789), .s(n9715), .op(
        n6149) );
  mux2_1 U11740 ( .ip1(\cache_data_B[1][84] ), .ip2(n9790), .s(n9715), .op(
        n6148) );
  mux2_1 U11741 ( .ip1(\cache_data_B[1][85] ), .ip2(n9791), .s(n9715), .op(
        n6147) );
  mux2_1 U11742 ( .ip1(\cache_data_B[1][86] ), .ip2(n9792), .s(n9715), .op(
        n6146) );
  mux2_1 U11743 ( .ip1(\cache_data_B[1][87] ), .ip2(n9794), .s(n9715), .op(
        n6145) );
  mux2_1 U11744 ( .ip1(\cache_data_B[1][88] ), .ip2(n9795), .s(n9716), .op(
        n6144) );
  mux2_1 U11745 ( .ip1(\cache_data_B[1][89] ), .ip2(n9796), .s(n9716), .op(
        n6143) );
  mux2_1 U11746 ( .ip1(\cache_data_B[1][90] ), .ip2(n9797), .s(n9716), .op(
        n6142) );
  mux2_1 U11747 ( .ip1(\cache_data_B[1][91] ), .ip2(n9798), .s(n9716), .op(
        n6141) );
  mux2_1 U11748 ( .ip1(\cache_data_B[1][92] ), .ip2(n9799), .s(n9716), .op(
        n6140) );
  mux2_1 U11749 ( .ip1(\cache_data_B[1][93] ), .ip2(n9800), .s(n9716), .op(
        n6139) );
  mux2_1 U11750 ( .ip1(\cache_data_B[1][94] ), .ip2(n9801), .s(n9716), .op(
        n6138) );
  mux2_1 U11751 ( .ip1(\cache_data_B[1][95] ), .ip2(n9803), .s(n9716), .op(
        n6137) );
  nand2_1 U11752 ( .ip1(n9717), .ip2(n9810), .op(n9718) );
  mux2_1 U11753 ( .ip1(n9770), .ip2(\cache_data_B[1][96] ), .s(n9718), .op(
        n6136) );
  mux2_1 U11754 ( .ip1(n9771), .ip2(\cache_data_B[1][97] ), .s(n9718), .op(
        n6135) );
  mux2_1 U11755 ( .ip1(n9772), .ip2(\cache_data_B[1][98] ), .s(n9718), .op(
        n6134) );
  mux2_1 U11756 ( .ip1(n9773), .ip2(\cache_data_B[1][99] ), .s(n9718), .op(
        n6133) );
  mux2_1 U11757 ( .ip1(n9774), .ip2(\cache_data_B[1][100] ), .s(n9718), .op(
        n6132) );
  mux2_1 U11758 ( .ip1(n9775), .ip2(\cache_data_B[1][101] ), .s(n9718), .op(
        n6131) );
  mux2_1 U11759 ( .ip1(n9776), .ip2(\cache_data_B[1][102] ), .s(n9718), .op(
        n6130) );
  mux2_1 U11760 ( .ip1(n9777), .ip2(\cache_data_B[1][103] ), .s(n9718), .op(
        n6129) );
  mux2_1 U11761 ( .ip1(n9778), .ip2(\cache_data_B[1][104] ), .s(n9718), .op(
        n6128) );
  mux2_1 U11762 ( .ip1(n9779), .ip2(\cache_data_B[1][105] ), .s(n9718), .op(
        n6127) );
  buf_1 U11763 ( .ip(n9718), .op(n9719) );
  mux2_1 U11764 ( .ip1(n9780), .ip2(\cache_data_B[1][106] ), .s(n9719), .op(
        n6126) );
  mux2_1 U11765 ( .ip1(n9781), .ip2(\cache_data_B[1][107] ), .s(n9718), .op(
        n6125) );
  mux2_1 U11766 ( .ip1(n9782), .ip2(\cache_data_B[1][108] ), .s(n9718), .op(
        n6124) );
  mux2_1 U11767 ( .ip1(n9783), .ip2(\cache_data_B[1][109] ), .s(n9718), .op(
        n6123) );
  mux2_1 U11768 ( .ip1(n9784), .ip2(\cache_data_B[1][110] ), .s(n9718), .op(
        n6122) );
  mux2_1 U11769 ( .ip1(n9785), .ip2(\cache_data_B[1][111] ), .s(n9718), .op(
        n6121) );
  mux2_1 U11770 ( .ip1(n9786), .ip2(\cache_data_B[1][112] ), .s(n9718), .op(
        n6120) );
  mux2_1 U11771 ( .ip1(n9787), .ip2(\cache_data_B[1][113] ), .s(n9718), .op(
        n6119) );
  mux2_1 U11772 ( .ip1(n9788), .ip2(\cache_data_B[1][114] ), .s(n9718), .op(
        n6118) );
  mux2_1 U11773 ( .ip1(n9789), .ip2(\cache_data_B[1][115] ), .s(n9718), .op(
        n6117) );
  mux2_1 U11774 ( .ip1(n9790), .ip2(\cache_data_B[1][116] ), .s(n9718), .op(
        n6116) );
  mux2_1 U11775 ( .ip1(n9791), .ip2(\cache_data_B[1][117] ), .s(n9718), .op(
        n6115) );
  mux2_1 U11776 ( .ip1(n9835), .ip2(\cache_data_B[1][118] ), .s(n9719), .op(
        n6114) );
  mux2_1 U11777 ( .ip1(n9794), .ip2(\cache_data_B[1][119] ), .s(n9719), .op(
        n6113) );
  mux2_1 U11778 ( .ip1(n9795), .ip2(\cache_data_B[1][120] ), .s(n9719), .op(
        n6112) );
  mux2_1 U11779 ( .ip1(n9796), .ip2(\cache_data_B[1][121] ), .s(n9719), .op(
        n6111) );
  mux2_1 U11780 ( .ip1(n9797), .ip2(\cache_data_B[1][122] ), .s(n9719), .op(
        n6110) );
  mux2_1 U11781 ( .ip1(n9798), .ip2(\cache_data_B[1][123] ), .s(n9719), .op(
        n6109) );
  mux2_1 U11782 ( .ip1(n9799), .ip2(\cache_data_B[1][124] ), .s(n9719), .op(
        n6108) );
  mux2_1 U11783 ( .ip1(n9800), .ip2(\cache_data_B[1][125] ), .s(n9719), .op(
        n6107) );
  mux2_1 U11784 ( .ip1(n9801), .ip2(\cache_data_B[1][126] ), .s(n9719), .op(
        n6106) );
  mux2_1 U11785 ( .ip1(n9803), .ip2(\cache_data_B[1][127] ), .s(n9719), .op(
        n6105) );
  nand2_1 U11786 ( .ip1(n9726), .ip2(n9756), .op(n9720) );
  mux2_1 U11787 ( .ip1(n9801), .ip2(\cache_data_B[2][30] ), .s(n9720), .op(
        n6104) );
  mux2_1 U11788 ( .ip1(n9803), .ip2(\cache_data_B[2][31] ), .s(n9720), .op(
        n6103) );
  mux2_1 U11789 ( .ip1(n9770), .ip2(\cache_data_B[2][0] ), .s(n9720), .op(
        n6102) );
  buf_1 U11790 ( .ip(n9720), .op(n9721) );
  mux2_1 U11791 ( .ip1(n9771), .ip2(\cache_data_B[2][1] ), .s(n9721), .op(
        n6101) );
  mux2_1 U11792 ( .ip1(n9772), .ip2(\cache_data_B[2][2] ), .s(n9720), .op(
        n6100) );
  mux2_1 U11793 ( .ip1(n9773), .ip2(\cache_data_B[2][3] ), .s(n9720), .op(
        n6099) );
  mux2_1 U11794 ( .ip1(n9774), .ip2(\cache_data_B[2][4] ), .s(n9720), .op(
        n6098) );
  mux2_1 U11795 ( .ip1(n9775), .ip2(\cache_data_B[2][5] ), .s(n9720), .op(
        n6097) );
  mux2_1 U11796 ( .ip1(n9776), .ip2(\cache_data_B[2][6] ), .s(n9720), .op(
        n6096) );
  mux2_1 U11797 ( .ip1(n9777), .ip2(\cache_data_B[2][7] ), .s(n9720), .op(
        n6095) );
  mux2_1 U11798 ( .ip1(n9778), .ip2(\cache_data_B[2][8] ), .s(n9720), .op(
        n6094) );
  mux2_1 U11799 ( .ip1(n9779), .ip2(\cache_data_B[2][9] ), .s(n9720), .op(
        n6093) );
  mux2_1 U11800 ( .ip1(n9780), .ip2(\cache_data_B[2][10] ), .s(n9720), .op(
        n6092) );
  mux2_1 U11801 ( .ip1(n9781), .ip2(\cache_data_B[2][11] ), .s(n9720), .op(
        n6091) );
  mux2_1 U11802 ( .ip1(n9782), .ip2(\cache_data_B[2][12] ), .s(n9721), .op(
        n6090) );
  mux2_1 U11803 ( .ip1(n9783), .ip2(\cache_data_B[2][13] ), .s(n9720), .op(
        n6089) );
  mux2_1 U11804 ( .ip1(n9784), .ip2(\cache_data_B[2][14] ), .s(n9720), .op(
        n6088) );
  mux2_1 U11805 ( .ip1(n9785), .ip2(\cache_data_B[2][15] ), .s(n9720), .op(
        n6087) );
  mux2_1 U11806 ( .ip1(n9786), .ip2(\cache_data_B[2][16] ), .s(n9720), .op(
        n6086) );
  mux2_1 U11807 ( .ip1(n9787), .ip2(\cache_data_B[2][17] ), .s(n9720), .op(
        n6085) );
  mux2_1 U11808 ( .ip1(n9788), .ip2(\cache_data_B[2][18] ), .s(n9721), .op(
        n6084) );
  mux2_1 U11809 ( .ip1(n9831), .ip2(\cache_data_B[2][19] ), .s(n9720), .op(
        n6083) );
  mux2_1 U11810 ( .ip1(n9790), .ip2(\cache_data_B[2][20] ), .s(n9721), .op(
        n6082) );
  mux2_1 U11811 ( .ip1(n9833), .ip2(\cache_data_B[2][21] ), .s(n9720), .op(
        n6081) );
  mux2_1 U11812 ( .ip1(n9835), .ip2(\cache_data_B[2][22] ), .s(n9720), .op(
        n6080) );
  mux2_1 U11813 ( .ip1(n9836), .ip2(\cache_data_B[2][23] ), .s(n9721), .op(
        n6079) );
  mux2_1 U11814 ( .ip1(n9837), .ip2(\cache_data_B[2][24] ), .s(n9721), .op(
        n6078) );
  mux2_1 U11815 ( .ip1(n9796), .ip2(\cache_data_B[2][25] ), .s(n9721), .op(
        n6077) );
  mux2_1 U11816 ( .ip1(n9797), .ip2(\cache_data_B[2][26] ), .s(n9721), .op(
        n6076) );
  mux2_1 U11817 ( .ip1(n9798), .ip2(\cache_data_B[2][27] ), .s(n9721), .op(
        n6075) );
  mux2_1 U11818 ( .ip1(n9799), .ip2(\cache_data_B[2][28] ), .s(n9721), .op(
        n6074) );
  mux2_1 U11819 ( .ip1(n9800), .ip2(\cache_data_B[2][29] ), .s(n9721), .op(
        n6073) );
  nand2_1 U11820 ( .ip1(n9726), .ip2(n9804), .op(n9722) );
  mux2_1 U11821 ( .ip1(n9770), .ip2(\cache_data_B[2][32] ), .s(n9722), .op(
        n6072) );
  mux2_1 U11822 ( .ip1(n9771), .ip2(\cache_data_B[2][33] ), .s(n9722), .op(
        n6071) );
  mux2_1 U11823 ( .ip1(n9772), .ip2(\cache_data_B[2][34] ), .s(n9722), .op(
        n6070) );
  mux2_1 U11824 ( .ip1(n9773), .ip2(\cache_data_B[2][35] ), .s(n9722), .op(
        n6069) );
  mux2_1 U11825 ( .ip1(n9774), .ip2(\cache_data_B[2][36] ), .s(n9722), .op(
        n6068) );
  mux2_1 U11826 ( .ip1(n9775), .ip2(\cache_data_B[2][37] ), .s(n9722), .op(
        n6067) );
  mux2_1 U11827 ( .ip1(n9776), .ip2(\cache_data_B[2][38] ), .s(n9722), .op(
        n6066) );
  mux2_1 U11828 ( .ip1(n9777), .ip2(\cache_data_B[2][39] ), .s(n9722), .op(
        n6065) );
  mux2_1 U11829 ( .ip1(n9778), .ip2(\cache_data_B[2][40] ), .s(n9722), .op(
        n6064) );
  buf_1 U11830 ( .ip(n9722), .op(n9723) );
  mux2_1 U11831 ( .ip1(n9779), .ip2(\cache_data_B[2][41] ), .s(n9723), .op(
        n6063) );
  mux2_1 U11832 ( .ip1(n9780), .ip2(\cache_data_B[2][42] ), .s(n9722), .op(
        n6062) );
  mux2_1 U11833 ( .ip1(n9781), .ip2(\cache_data_B[2][43] ), .s(n9722), .op(
        n6061) );
  mux2_1 U11834 ( .ip1(n9782), .ip2(\cache_data_B[2][44] ), .s(n9722), .op(
        n6060) );
  mux2_1 U11835 ( .ip1(n9783), .ip2(\cache_data_B[2][45] ), .s(n9722), .op(
        n6059) );
  mux2_1 U11836 ( .ip1(n9784), .ip2(\cache_data_B[2][46] ), .s(n9722), .op(
        n6058) );
  mux2_1 U11837 ( .ip1(n9785), .ip2(\cache_data_B[2][47] ), .s(n9722), .op(
        n6057) );
  mux2_1 U11838 ( .ip1(n9786), .ip2(\cache_data_B[2][48] ), .s(n9722), .op(
        n6056) );
  mux2_1 U11839 ( .ip1(n9787), .ip2(\cache_data_B[2][49] ), .s(n9723), .op(
        n6055) );
  mux2_1 U11840 ( .ip1(n9788), .ip2(\cache_data_B[2][50] ), .s(n9722), .op(
        n6054) );
  mux2_1 U11841 ( .ip1(n9789), .ip2(\cache_data_B[2][51] ), .s(n9722), .op(
        n6053) );
  mux2_1 U11842 ( .ip1(n9832), .ip2(\cache_data_B[2][52] ), .s(n9723), .op(
        n6052) );
  mux2_1 U11843 ( .ip1(n9833), .ip2(\cache_data_B[2][53] ), .s(n9722), .op(
        n6051) );
  mux2_1 U11844 ( .ip1(n9792), .ip2(\cache_data_B[2][54] ), .s(n9722), .op(
        n6050) );
  mux2_1 U11845 ( .ip1(n9836), .ip2(\cache_data_B[2][55] ), .s(n9722), .op(
        n6049) );
  mux2_1 U11846 ( .ip1(n9837), .ip2(\cache_data_B[2][56] ), .s(n9723), .op(
        n6048) );
  mux2_1 U11847 ( .ip1(n9796), .ip2(\cache_data_B[2][57] ), .s(n9723), .op(
        n6047) );
  mux2_1 U11848 ( .ip1(n9797), .ip2(\cache_data_B[2][58] ), .s(n9723), .op(
        n6046) );
  mux2_1 U11849 ( .ip1(n9798), .ip2(\cache_data_B[2][59] ), .s(n9723), .op(
        n6045) );
  mux2_1 U11850 ( .ip1(n9799), .ip2(\cache_data_B[2][60] ), .s(n9723), .op(
        n6044) );
  mux2_1 U11851 ( .ip1(n9800), .ip2(\cache_data_B[2][61] ), .s(n9723), .op(
        n6043) );
  mux2_1 U11852 ( .ip1(n9801), .ip2(\cache_data_B[2][62] ), .s(n9723), .op(
        n6042) );
  mux2_1 U11853 ( .ip1(n9803), .ip2(\cache_data_B[2][63] ), .s(n9723), .op(
        n6041) );
  nor2_1 U11854 ( .ip1(n9864), .ip2(n9761), .op(n9724) );
  buf_1 U11855 ( .ip(n9724), .op(n9725) );
  mux2_1 U11856 ( .ip1(\cache_data_B[2][64] ), .ip2(n9770), .s(n9725), .op(
        n6040) );
  mux2_1 U11857 ( .ip1(\cache_data_B[2][65] ), .ip2(n9771), .s(n9724), .op(
        n6039) );
  mux2_1 U11858 ( .ip1(\cache_data_B[2][66] ), .ip2(n9772), .s(n9724), .op(
        n6038) );
  mux2_1 U11859 ( .ip1(\cache_data_B[2][67] ), .ip2(n9773), .s(n9724), .op(
        n6037) );
  mux2_1 U11860 ( .ip1(\cache_data_B[2][68] ), .ip2(n9774), .s(n9724), .op(
        n6036) );
  mux2_1 U11861 ( .ip1(\cache_data_B[2][69] ), .ip2(n9775), .s(n9724), .op(
        n6035) );
  mux2_1 U11862 ( .ip1(\cache_data_B[2][70] ), .ip2(n9776), .s(n9724), .op(
        n6034) );
  mux2_1 U11863 ( .ip1(\cache_data_B[2][71] ), .ip2(n9777), .s(n9724), .op(
        n6033) );
  mux2_1 U11864 ( .ip1(\cache_data_B[2][72] ), .ip2(n9778), .s(n9724), .op(
        n6032) );
  mux2_1 U11865 ( .ip1(\cache_data_B[2][73] ), .ip2(n9779), .s(n9725), .op(
        n6031) );
  mux2_1 U11866 ( .ip1(\cache_data_B[2][74] ), .ip2(n9780), .s(n9725), .op(
        n6030) );
  mux2_1 U11867 ( .ip1(\cache_data_B[2][75] ), .ip2(n9781), .s(n9724), .op(
        n6029) );
  mux2_1 U11868 ( .ip1(\cache_data_B[2][76] ), .ip2(n9782), .s(n9724), .op(
        n6028) );
  mux2_1 U11869 ( .ip1(\cache_data_B[2][77] ), .ip2(n9783), .s(n9724), .op(
        n6027) );
  mux2_1 U11870 ( .ip1(\cache_data_B[2][78] ), .ip2(n9784), .s(n9724), .op(
        n6026) );
  mux2_1 U11871 ( .ip1(\cache_data_B[2][79] ), .ip2(n9785), .s(n9724), .op(
        n6025) );
  mux2_1 U11872 ( .ip1(\cache_data_B[2][80] ), .ip2(n9786), .s(n9724), .op(
        n6024) );
  mux2_1 U11873 ( .ip1(\cache_data_B[2][81] ), .ip2(n9787), .s(n9724), .op(
        n6023) );
  mux2_1 U11874 ( .ip1(\cache_data_B[2][82] ), .ip2(n9788), .s(n9724), .op(
        n6022) );
  mux2_1 U11875 ( .ip1(\cache_data_B[2][83] ), .ip2(n9831), .s(n9724), .op(
        n6021) );
  mux2_1 U11876 ( .ip1(\cache_data_B[2][84] ), .ip2(n9832), .s(n9724), .op(
        n6020) );
  mux2_1 U11877 ( .ip1(\cache_data_B[2][85] ), .ip2(n9833), .s(n9724), .op(
        n6019) );
  mux2_1 U11878 ( .ip1(\cache_data_B[2][86] ), .ip2(n9835), .s(n9724), .op(
        n6018) );
  mux2_1 U11879 ( .ip1(\cache_data_B[2][87] ), .ip2(n9836), .s(n9724), .op(
        n6017) );
  mux2_1 U11880 ( .ip1(\cache_data_B[2][88] ), .ip2(n9837), .s(n9725), .op(
        n6016) );
  mux2_1 U11881 ( .ip1(\cache_data_B[2][89] ), .ip2(n9796), .s(n9725), .op(
        n6015) );
  mux2_1 U11882 ( .ip1(\cache_data_B[2][90] ), .ip2(n9797), .s(n9725), .op(
        n6014) );
  mux2_1 U11883 ( .ip1(\cache_data_B[2][91] ), .ip2(n9798), .s(n9725), .op(
        n6013) );
  mux2_1 U11884 ( .ip1(\cache_data_B[2][92] ), .ip2(n9799), .s(n9725), .op(
        n6012) );
  mux2_1 U11885 ( .ip1(\cache_data_B[2][93] ), .ip2(n9800), .s(n9725), .op(
        n6011) );
  mux2_1 U11886 ( .ip1(\cache_data_B[2][94] ), .ip2(n9801), .s(n9725), .op(
        n6010) );
  mux2_1 U11887 ( .ip1(\cache_data_B[2][95] ), .ip2(n9803), .s(n9725), .op(
        n6009) );
  nand2_1 U11888 ( .ip1(n9726), .ip2(n9810), .op(n9727) );
  mux2_1 U11889 ( .ip1(n9770), .ip2(\cache_data_B[2][96] ), .s(n9727), .op(
        n6008) );
  mux2_1 U11890 ( .ip1(n9771), .ip2(\cache_data_B[2][97] ), .s(n9727), .op(
        n6007) );
  mux2_1 U11891 ( .ip1(n9772), .ip2(\cache_data_B[2][98] ), .s(n9727), .op(
        n6006) );
  mux2_1 U11892 ( .ip1(n9773), .ip2(\cache_data_B[2][99] ), .s(n9727), .op(
        n6005) );
  buf_1 U11893 ( .ip(n9727), .op(n9728) );
  mux2_1 U11894 ( .ip1(n9774), .ip2(\cache_data_B[2][100] ), .s(n9728), .op(
        n6004) );
  mux2_1 U11895 ( .ip1(n9775), .ip2(\cache_data_B[2][101] ), .s(n9727), .op(
        n6003) );
  mux2_1 U11896 ( .ip1(n9776), .ip2(\cache_data_B[2][102] ), .s(n9727), .op(
        n6002) );
  mux2_1 U11897 ( .ip1(n9777), .ip2(\cache_data_B[2][103] ), .s(n9727), .op(
        n6001) );
  mux2_1 U11898 ( .ip1(n9778), .ip2(\cache_data_B[2][104] ), .s(n9727), .op(
        n6000) );
  mux2_1 U11899 ( .ip1(n9779), .ip2(\cache_data_B[2][105] ), .s(n9727), .op(
        n5999) );
  mux2_1 U11900 ( .ip1(n9780), .ip2(\cache_data_B[2][106] ), .s(n9727), .op(
        n5998) );
  mux2_1 U11901 ( .ip1(n9781), .ip2(\cache_data_B[2][107] ), .s(n9727), .op(
        n5997) );
  mux2_1 U11902 ( .ip1(n9782), .ip2(\cache_data_B[2][108] ), .s(n9727), .op(
        n5996) );
  mux2_1 U11903 ( .ip1(n9783), .ip2(\cache_data_B[2][109] ), .s(n9727), .op(
        n5995) );
  mux2_1 U11904 ( .ip1(n9784), .ip2(\cache_data_B[2][110] ), .s(n9727), .op(
        n5994) );
  mux2_1 U11905 ( .ip1(n9785), .ip2(\cache_data_B[2][111] ), .s(n9727), .op(
        n5993) );
  mux2_1 U11906 ( .ip1(n9786), .ip2(\cache_data_B[2][112] ), .s(n9727), .op(
        n5992) );
  mux2_1 U11907 ( .ip1(n9787), .ip2(\cache_data_B[2][113] ), .s(n9727), .op(
        n5991) );
  mux2_1 U11908 ( .ip1(n9788), .ip2(\cache_data_B[2][114] ), .s(n9727), .op(
        n5990) );
  mux2_1 U11909 ( .ip1(n9831), .ip2(\cache_data_B[2][115] ), .s(n9728), .op(
        n5989) );
  mux2_1 U11910 ( .ip1(n9832), .ip2(\cache_data_B[2][116] ), .s(n9728), .op(
        n5988) );
  mux2_1 U11911 ( .ip1(n9833), .ip2(\cache_data_B[2][117] ), .s(n9728), .op(
        n5987) );
  mux2_1 U11912 ( .ip1(n9835), .ip2(\cache_data_B[2][118] ), .s(n9728), .op(
        n5986) );
  mux2_1 U11913 ( .ip1(n9794), .ip2(\cache_data_B[2][119] ), .s(n9727), .op(
        n5985) );
  mux2_1 U11914 ( .ip1(n9795), .ip2(\cache_data_B[2][120] ), .s(n9727), .op(
        n5984) );
  mux2_1 U11915 ( .ip1(n9796), .ip2(\cache_data_B[2][121] ), .s(n9727), .op(
        n5983) );
  mux2_1 U11916 ( .ip1(n9797), .ip2(\cache_data_B[2][122] ), .s(n9728), .op(
        n5982) );
  mux2_1 U11917 ( .ip1(n9798), .ip2(\cache_data_B[2][123] ), .s(n9728), .op(
        n5981) );
  mux2_1 U11918 ( .ip1(n9799), .ip2(\cache_data_B[2][124] ), .s(n9728), .op(
        n5980) );
  mux2_1 U11919 ( .ip1(n9800), .ip2(\cache_data_B[2][125] ), .s(n9728), .op(
        n5979) );
  mux2_1 U11920 ( .ip1(n9801), .ip2(\cache_data_B[2][126] ), .s(n9728), .op(
        n5978) );
  mux2_1 U11921 ( .ip1(n9803), .ip2(\cache_data_B[2][127] ), .s(n9728), .op(
        n5977) );
  nand2_1 U11922 ( .ip1(n9735), .ip2(n9756), .op(n9729) );
  mux2_1 U11923 ( .ip1(n9771), .ip2(\cache_data_B[3][1] ), .s(n9729), .op(
        n5976) );
  mux2_1 U11924 ( .ip1(n9772), .ip2(\cache_data_B[3][2] ), .s(n9729), .op(
        n5975) );
  mux2_1 U11925 ( .ip1(n9773), .ip2(\cache_data_B[3][3] ), .s(n9729), .op(
        n5974) );
  mux2_1 U11926 ( .ip1(n9774), .ip2(\cache_data_B[3][4] ), .s(n9729), .op(
        n5973) );
  mux2_1 U11927 ( .ip1(n9775), .ip2(\cache_data_B[3][5] ), .s(n9729), .op(
        n5972) );
  mux2_1 U11928 ( .ip1(n9776), .ip2(\cache_data_B[3][6] ), .s(n9729), .op(
        n5971) );
  mux2_1 U11929 ( .ip1(n9777), .ip2(\cache_data_B[3][7] ), .s(n9729), .op(
        n5970) );
  mux2_1 U11930 ( .ip1(n9778), .ip2(\cache_data_B[3][8] ), .s(n9729), .op(
        n5969) );
  mux2_1 U11931 ( .ip1(n9779), .ip2(\cache_data_B[3][9] ), .s(n9729), .op(
        n5968) );
  buf_1 U11932 ( .ip(n9729), .op(n9730) );
  mux2_1 U11933 ( .ip1(n9780), .ip2(\cache_data_B[3][10] ), .s(n9730), .op(
        n5967) );
  mux2_1 U11934 ( .ip1(n9781), .ip2(\cache_data_B[3][11] ), .s(n9729), .op(
        n5966) );
  mux2_1 U11935 ( .ip1(n9782), .ip2(\cache_data_B[3][12] ), .s(n9729), .op(
        n5965) );
  mux2_1 U11936 ( .ip1(n9783), .ip2(\cache_data_B[3][13] ), .s(n9729), .op(
        n5964) );
  mux2_1 U11937 ( .ip1(n9784), .ip2(\cache_data_B[3][14] ), .s(n9729), .op(
        n5963) );
  mux2_1 U11938 ( .ip1(n9785), .ip2(\cache_data_B[3][15] ), .s(n9730), .op(
        n5962) );
  mux2_1 U11939 ( .ip1(n9786), .ip2(\cache_data_B[3][16] ), .s(n9729), .op(
        n5961) );
  mux2_1 U11940 ( .ip1(n9787), .ip2(\cache_data_B[3][17] ), .s(n9729), .op(
        n5960) );
  mux2_1 U11941 ( .ip1(n9788), .ip2(\cache_data_B[3][18] ), .s(n9729), .op(
        n5959) );
  mux2_1 U11942 ( .ip1(n9831), .ip2(\cache_data_B[3][19] ), .s(n9729), .op(
        n5958) );
  mux2_1 U11943 ( .ip1(n9832), .ip2(\cache_data_B[3][20] ), .s(n9729), .op(
        n5957) );
  mux2_1 U11944 ( .ip1(n9791), .ip2(\cache_data_B[3][21] ), .s(n9729), .op(
        n5956) );
  mux2_1 U11945 ( .ip1(n9792), .ip2(\cache_data_B[3][22] ), .s(n9729), .op(
        n5955) );
  mux2_1 U11946 ( .ip1(n9794), .ip2(\cache_data_B[3][23] ), .s(n9729), .op(
        n5954) );
  mux2_1 U11947 ( .ip1(n9795), .ip2(\cache_data_B[3][24] ), .s(n9730), .op(
        n5953) );
  mux2_1 U11948 ( .ip1(n9796), .ip2(\cache_data_B[3][25] ), .s(n9730), .op(
        n5952) );
  mux2_1 U11949 ( .ip1(n9797), .ip2(\cache_data_B[3][26] ), .s(n9730), .op(
        n5951) );
  mux2_1 U11950 ( .ip1(n9798), .ip2(\cache_data_B[3][27] ), .s(n9730), .op(
        n5950) );
  mux2_1 U11951 ( .ip1(n9799), .ip2(\cache_data_B[3][28] ), .s(n9730), .op(
        n5949) );
  mux2_1 U11952 ( .ip1(n9800), .ip2(\cache_data_B[3][29] ), .s(n9730), .op(
        n5948) );
  mux2_1 U11953 ( .ip1(n9801), .ip2(\cache_data_B[3][30] ), .s(n9730), .op(
        n5947) );
  mux2_1 U11954 ( .ip1(n9803), .ip2(\cache_data_B[3][31] ), .s(n9730), .op(
        n5946) );
  mux2_1 U11955 ( .ip1(n9770), .ip2(\cache_data_B[3][0] ), .s(n9730), .op(
        n5945) );
  nand2_1 U11956 ( .ip1(n9735), .ip2(n9804), .op(n9731) );
  mux2_1 U11957 ( .ip1(n9770), .ip2(\cache_data_B[3][32] ), .s(n9731), .op(
        n5944) );
  mux2_1 U11958 ( .ip1(n9771), .ip2(\cache_data_B[3][33] ), .s(n9731), .op(
        n5943) );
  mux2_1 U11959 ( .ip1(n9772), .ip2(\cache_data_B[3][34] ), .s(n9731), .op(
        n5942) );
  mux2_1 U11960 ( .ip1(n9773), .ip2(\cache_data_B[3][35] ), .s(n9731), .op(
        n5941) );
  mux2_1 U11961 ( .ip1(n9774), .ip2(\cache_data_B[3][36] ), .s(n9731), .op(
        n5940) );
  mux2_1 U11962 ( .ip1(n9775), .ip2(\cache_data_B[3][37] ), .s(n9731), .op(
        n5939) );
  mux2_1 U11963 ( .ip1(n9776), .ip2(\cache_data_B[3][38] ), .s(n9731), .op(
        n5938) );
  mux2_1 U11964 ( .ip1(n9777), .ip2(\cache_data_B[3][39] ), .s(n9731), .op(
        n5937) );
  mux2_1 U11965 ( .ip1(n9778), .ip2(\cache_data_B[3][40] ), .s(n9731), .op(
        n5936) );
  mux2_1 U11966 ( .ip1(n9779), .ip2(\cache_data_B[3][41] ), .s(n9731), .op(
        n5935) );
  buf_1 U11967 ( .ip(n9731), .op(n9732) );
  mux2_1 U11968 ( .ip1(n9780), .ip2(\cache_data_B[3][42] ), .s(n9732), .op(
        n5934) );
  mux2_1 U11969 ( .ip1(n9781), .ip2(\cache_data_B[3][43] ), .s(n9731), .op(
        n5933) );
  mux2_1 U11970 ( .ip1(n9782), .ip2(\cache_data_B[3][44] ), .s(n9731), .op(
        n5932) );
  mux2_1 U11971 ( .ip1(n9783), .ip2(\cache_data_B[3][45] ), .s(n9732), .op(
        n5931) );
  mux2_1 U11972 ( .ip1(n9784), .ip2(\cache_data_B[3][46] ), .s(n9732), .op(
        n5930) );
  mux2_1 U11973 ( .ip1(n9785), .ip2(\cache_data_B[3][47] ), .s(n9731), .op(
        n5929) );
  mux2_1 U11974 ( .ip1(n9786), .ip2(\cache_data_B[3][48] ), .s(n9731), .op(
        n5928) );
  mux2_1 U11975 ( .ip1(n9787), .ip2(\cache_data_B[3][49] ), .s(n9731), .op(
        n5927) );
  mux2_1 U11976 ( .ip1(n9788), .ip2(\cache_data_B[3][50] ), .s(n9731), .op(
        n5926) );
  mux2_1 U11977 ( .ip1(n9789), .ip2(\cache_data_B[3][51] ), .s(n9731), .op(
        n5925) );
  mux2_1 U11978 ( .ip1(n9832), .ip2(\cache_data_B[3][52] ), .s(n9731), .op(
        n5924) );
  mux2_1 U11979 ( .ip1(n9791), .ip2(\cache_data_B[3][53] ), .s(n9731), .op(
        n5923) );
  mux2_1 U11980 ( .ip1(n9792), .ip2(\cache_data_B[3][54] ), .s(n9732), .op(
        n5922) );
  mux2_1 U11981 ( .ip1(n9794), .ip2(\cache_data_B[3][55] ), .s(n9732), .op(
        n5921) );
  mux2_1 U11982 ( .ip1(n9837), .ip2(\cache_data_B[3][56] ), .s(n9731), .op(
        n5920) );
  mux2_1 U11983 ( .ip1(n9796), .ip2(\cache_data_B[3][57] ), .s(n9731), .op(
        n5919) );
  mux2_1 U11984 ( .ip1(n9797), .ip2(\cache_data_B[3][58] ), .s(n9732), .op(
        n5918) );
  mux2_1 U11985 ( .ip1(n9798), .ip2(\cache_data_B[3][59] ), .s(n9732), .op(
        n5917) );
  mux2_1 U11986 ( .ip1(n9799), .ip2(\cache_data_B[3][60] ), .s(n9732), .op(
        n5916) );
  mux2_1 U11987 ( .ip1(n9800), .ip2(\cache_data_B[3][61] ), .s(n9732), .op(
        n5915) );
  mux2_1 U11988 ( .ip1(n9801), .ip2(\cache_data_B[3][62] ), .s(n9732), .op(
        n5914) );
  mux2_1 U11989 ( .ip1(n9803), .ip2(\cache_data_B[3][63] ), .s(n9732), .op(
        n5913) );
  nor2_1 U11990 ( .ip1(n9866), .ip2(n9761), .op(n9733) );
  buf_1 U11991 ( .ip(n9733), .op(n9734) );
  mux2_1 U11992 ( .ip1(\cache_data_B[3][64] ), .ip2(n9812), .s(n9734), .op(
        n5912) );
  mux2_1 U11993 ( .ip1(\cache_data_B[3][65] ), .ip2(n9771), .s(n9733), .op(
        n5911) );
  mux2_1 U11994 ( .ip1(\cache_data_B[3][66] ), .ip2(n9772), .s(n9733), .op(
        n5910) );
  mux2_1 U11995 ( .ip1(\cache_data_B[3][67] ), .ip2(n9773), .s(n9733), .op(
        n5909) );
  mux2_1 U11996 ( .ip1(\cache_data_B[3][68] ), .ip2(n9774), .s(n9733), .op(
        n5908) );
  mux2_1 U11997 ( .ip1(\cache_data_B[3][69] ), .ip2(n9775), .s(n9733), .op(
        n5907) );
  mux2_1 U11998 ( .ip1(\cache_data_B[3][70] ), .ip2(n9776), .s(n9733), .op(
        n5906) );
  mux2_1 U11999 ( .ip1(\cache_data_B[3][71] ), .ip2(n9777), .s(n9733), .op(
        n5905) );
  mux2_1 U12000 ( .ip1(\cache_data_B[3][72] ), .ip2(n9778), .s(n9733), .op(
        n5904) );
  mux2_1 U12001 ( .ip1(\cache_data_B[3][73] ), .ip2(n9779), .s(n9734), .op(
        n5903) );
  mux2_1 U12002 ( .ip1(\cache_data_B[3][74] ), .ip2(n9780), .s(n9734), .op(
        n5902) );
  mux2_1 U12003 ( .ip1(\cache_data_B[3][75] ), .ip2(n9781), .s(n9733), .op(
        n5901) );
  mux2_1 U12004 ( .ip1(\cache_data_B[3][76] ), .ip2(n9782), .s(n9733), .op(
        n5900) );
  mux2_1 U12005 ( .ip1(\cache_data_B[3][77] ), .ip2(n9783), .s(n9733), .op(
        n5899) );
  mux2_1 U12006 ( .ip1(\cache_data_B[3][78] ), .ip2(n9784), .s(n9733), .op(
        n5898) );
  mux2_1 U12007 ( .ip1(\cache_data_B[3][79] ), .ip2(n9785), .s(n9733), .op(
        n5897) );
  mux2_1 U12008 ( .ip1(\cache_data_B[3][80] ), .ip2(n9786), .s(n9733), .op(
        n5896) );
  mux2_1 U12009 ( .ip1(\cache_data_B[3][81] ), .ip2(n9829), .s(n9733), .op(
        n5895) );
  mux2_1 U12010 ( .ip1(\cache_data_B[3][82] ), .ip2(n9830), .s(n9733), .op(
        n5894) );
  mux2_1 U12011 ( .ip1(\cache_data_B[3][83] ), .ip2(n9831), .s(n9733), .op(
        n5893) );
  mux2_1 U12012 ( .ip1(\cache_data_B[3][84] ), .ip2(n9790), .s(n9733), .op(
        n5892) );
  mux2_1 U12013 ( .ip1(\cache_data_B[3][85] ), .ip2(n9791), .s(n9733), .op(
        n5891) );
  mux2_1 U12014 ( .ip1(\cache_data_B[3][86] ), .ip2(n9792), .s(n9733), .op(
        n5890) );
  mux2_1 U12015 ( .ip1(\cache_data_B[3][87] ), .ip2(n9794), .s(n9733), .op(
        n5889) );
  mux2_1 U12016 ( .ip1(\cache_data_B[3][88] ), .ip2(n9795), .s(n9734), .op(
        n5888) );
  mux2_1 U12017 ( .ip1(\cache_data_B[3][89] ), .ip2(n9838), .s(n9734), .op(
        n5887) );
  mux2_1 U12018 ( .ip1(\cache_data_B[3][90] ), .ip2(n9839), .s(n9734), .op(
        n5886) );
  mux2_1 U12019 ( .ip1(\cache_data_B[3][91] ), .ip2(n9840), .s(n9734), .op(
        n5885) );
  mux2_1 U12020 ( .ip1(\cache_data_B[3][92] ), .ip2(n9841), .s(n9734), .op(
        n5884) );
  mux2_1 U12021 ( .ip1(\cache_data_B[3][93] ), .ip2(n9842), .s(n9734), .op(
        n5883) );
  mux2_1 U12022 ( .ip1(\cache_data_B[3][94] ), .ip2(n9843), .s(n9734), .op(
        n5882) );
  mux2_1 U12023 ( .ip1(\cache_data_B[3][95] ), .ip2(n9845), .s(n9734), .op(
        n5881) );
  nand2_1 U12024 ( .ip1(n9735), .ip2(n9810), .op(n9736) );
  mux2_1 U12025 ( .ip1(n9816), .ip2(\cache_data_B[3][100] ), .s(n9736), .op(
        n5880) );
  mux2_1 U12026 ( .ip1(n9817), .ip2(\cache_data_B[3][101] ), .s(n9736), .op(
        n5879) );
  mux2_1 U12027 ( .ip1(n9818), .ip2(\cache_data_B[3][102] ), .s(n9736), .op(
        n5878) );
  mux2_1 U12028 ( .ip1(n9819), .ip2(\cache_data_B[3][103] ), .s(n9736), .op(
        n5877) );
  mux2_1 U12029 ( .ip1(n9820), .ip2(\cache_data_B[3][104] ), .s(n9736), .op(
        n5876) );
  mux2_1 U12030 ( .ip1(n9821), .ip2(\cache_data_B[3][105] ), .s(n9736), .op(
        n5875) );
  mux2_1 U12031 ( .ip1(n9822), .ip2(\cache_data_B[3][106] ), .s(n9736), .op(
        n5874) );
  mux2_1 U12032 ( .ip1(n9823), .ip2(\cache_data_B[3][107] ), .s(n9736), .op(
        n5873) );
  mux2_1 U12033 ( .ip1(n9824), .ip2(\cache_data_B[3][108] ), .s(n9736), .op(
        n5872) );
  mux2_1 U12034 ( .ip1(n9825), .ip2(\cache_data_B[3][109] ), .s(n9736), .op(
        n5871) );
  buf_1 U12035 ( .ip(n9736), .op(n9737) );
  mux2_1 U12036 ( .ip1(n9826), .ip2(\cache_data_B[3][110] ), .s(n9737), .op(
        n5870) );
  mux2_1 U12037 ( .ip1(n9827), .ip2(\cache_data_B[3][111] ), .s(n9736), .op(
        n5869) );
  mux2_1 U12038 ( .ip1(n9828), .ip2(\cache_data_B[3][112] ), .s(n9736), .op(
        n5868) );
  mux2_1 U12039 ( .ip1(n9829), .ip2(\cache_data_B[3][113] ), .s(n9736), .op(
        n5867) );
  mux2_1 U12040 ( .ip1(n9830), .ip2(\cache_data_B[3][114] ), .s(n9737), .op(
        n5866) );
  mux2_1 U12041 ( .ip1(n9831), .ip2(\cache_data_B[3][115] ), .s(n9736), .op(
        n5865) );
  mux2_1 U12042 ( .ip1(n9832), .ip2(\cache_data_B[3][116] ), .s(n9736), .op(
        n5864) );
  mux2_1 U12043 ( .ip1(n9833), .ip2(\cache_data_B[3][117] ), .s(n9736), .op(
        n5863) );
  mux2_1 U12044 ( .ip1(n9835), .ip2(\cache_data_B[3][118] ), .s(n9736), .op(
        n5862) );
  mux2_1 U12045 ( .ip1(n9836), .ip2(\cache_data_B[3][119] ), .s(n9736), .op(
        n5861) );
  mux2_1 U12046 ( .ip1(n9837), .ip2(\cache_data_B[3][120] ), .s(n9736), .op(
        n5860) );
  mux2_1 U12047 ( .ip1(n9838), .ip2(\cache_data_B[3][121] ), .s(n9737), .op(
        n5859) );
  mux2_1 U12048 ( .ip1(n9839), .ip2(\cache_data_B[3][122] ), .s(n9736), .op(
        n5858) );
  mux2_1 U12049 ( .ip1(n9840), .ip2(\cache_data_B[3][123] ), .s(n9736), .op(
        n5857) );
  mux2_1 U12050 ( .ip1(n9841), .ip2(\cache_data_B[3][124] ), .s(n9737), .op(
        n5856) );
  mux2_1 U12051 ( .ip1(n9842), .ip2(\cache_data_B[3][125] ), .s(n9737), .op(
        n5855) );
  mux2_1 U12052 ( .ip1(n9843), .ip2(\cache_data_B[3][126] ), .s(n9737), .op(
        n5854) );
  mux2_1 U12053 ( .ip1(n9845), .ip2(\cache_data_B[3][127] ), .s(n9737), .op(
        n5853) );
  mux2_1 U12054 ( .ip1(n9812), .ip2(\cache_data_B[3][96] ), .s(n9737), .op(
        n5852) );
  mux2_1 U12055 ( .ip1(n9813), .ip2(\cache_data_B[3][97] ), .s(n9737), .op(
        n5851) );
  mux2_1 U12056 ( .ip1(n9814), .ip2(\cache_data_B[3][98] ), .s(n9737), .op(
        n5850) );
  mux2_1 U12057 ( .ip1(n9815), .ip2(\cache_data_B[3][99] ), .s(n9737), .op(
        n5849) );
  nor2_1 U12058 ( .ip1(n9868), .ip2(n9768), .op(n9738) );
  buf_1 U12059 ( .ip(n9738), .op(n9739) );
  mux2_1 U12060 ( .ip1(\cache_data_B[4][0] ), .ip2(n9812), .s(n9739), .op(
        n5848) );
  mux2_1 U12061 ( .ip1(\cache_data_B[4][1] ), .ip2(n9813), .s(n9738), .op(
        n5847) );
  mux2_1 U12062 ( .ip1(\cache_data_B[4][2] ), .ip2(n9814), .s(n9738), .op(
        n5846) );
  mux2_1 U12063 ( .ip1(\cache_data_B[4][3] ), .ip2(n9815), .s(n9738), .op(
        n5845) );
  mux2_1 U12064 ( .ip1(\cache_data_B[4][4] ), .ip2(n9816), .s(n9738), .op(
        n5844) );
  mux2_1 U12065 ( .ip1(\cache_data_B[4][5] ), .ip2(n9817), .s(n9738), .op(
        n5843) );
  mux2_1 U12066 ( .ip1(\cache_data_B[4][6] ), .ip2(n9818), .s(n9738), .op(
        n5842) );
  mux2_1 U12067 ( .ip1(\cache_data_B[4][7] ), .ip2(n9819), .s(n9738), .op(
        n5841) );
  mux2_1 U12068 ( .ip1(\cache_data_B[4][8] ), .ip2(n9820), .s(n9738), .op(
        n5840) );
  mux2_1 U12069 ( .ip1(\cache_data_B[4][9] ), .ip2(n9821), .s(n9739), .op(
        n5839) );
  mux2_1 U12070 ( .ip1(\cache_data_B[4][10] ), .ip2(n9822), .s(n9739), .op(
        n5838) );
  mux2_1 U12071 ( .ip1(\cache_data_B[4][11] ), .ip2(n9823), .s(n9738), .op(
        n5837) );
  mux2_1 U12072 ( .ip1(\cache_data_B[4][12] ), .ip2(n9824), .s(n9738), .op(
        n5836) );
  mux2_1 U12073 ( .ip1(\cache_data_B[4][13] ), .ip2(n9825), .s(n9738), .op(
        n5835) );
  mux2_1 U12074 ( .ip1(\cache_data_B[4][14] ), .ip2(n9826), .s(n9738), .op(
        n5834) );
  mux2_1 U12075 ( .ip1(\cache_data_B[4][15] ), .ip2(n9827), .s(n9738), .op(
        n5833) );
  mux2_1 U12076 ( .ip1(\cache_data_B[4][16] ), .ip2(n9828), .s(n9738), .op(
        n5832) );
  mux2_1 U12077 ( .ip1(\cache_data_B[4][17] ), .ip2(n9829), .s(n9738), .op(
        n5831) );
  mux2_1 U12078 ( .ip1(\cache_data_B[4][18] ), .ip2(n9830), .s(n9738), .op(
        n5830) );
  mux2_1 U12079 ( .ip1(\cache_data_B[4][19] ), .ip2(n9831), .s(n9738), .op(
        n5829) );
  mux2_1 U12080 ( .ip1(\cache_data_B[4][20] ), .ip2(n9790), .s(n9738), .op(
        n5828) );
  mux2_1 U12081 ( .ip1(\cache_data_B[4][21] ), .ip2(n9791), .s(n9738), .op(
        n5827) );
  mux2_1 U12082 ( .ip1(\cache_data_B[4][22] ), .ip2(n9792), .s(n9738), .op(
        n5826) );
  mux2_1 U12083 ( .ip1(\cache_data_B[4][23] ), .ip2(n9794), .s(n9738), .op(
        n5825) );
  mux2_1 U12084 ( .ip1(\cache_data_B[4][24] ), .ip2(n9795), .s(n9739), .op(
        n5824) );
  mux2_1 U12085 ( .ip1(\cache_data_B[4][25] ), .ip2(n9838), .s(n9739), .op(
        n5823) );
  mux2_1 U12086 ( .ip1(\cache_data_B[4][26] ), .ip2(n9839), .s(n9739), .op(
        n5822) );
  mux2_1 U12087 ( .ip1(\cache_data_B[4][27] ), .ip2(n9840), .s(n9739), .op(
        n5821) );
  mux2_1 U12088 ( .ip1(\cache_data_B[4][28] ), .ip2(n9841), .s(n9739), .op(
        n5820) );
  mux2_1 U12089 ( .ip1(\cache_data_B[4][29] ), .ip2(n9842), .s(n9739), .op(
        n5819) );
  mux2_1 U12090 ( .ip1(\cache_data_B[4][30] ), .ip2(n9843), .s(n9739), .op(
        n5818) );
  mux2_1 U12091 ( .ip1(\cache_data_B[4][31] ), .ip2(n9845), .s(n9739), .op(
        n5817) );
  nand2_1 U12092 ( .ip1(n9744), .ip2(n9804), .op(n9740) );
  mux2_1 U12093 ( .ip1(n9812), .ip2(\cache_data_B[4][32] ), .s(n9740), .op(
        n5816) );
  mux2_1 U12094 ( .ip1(n9813), .ip2(\cache_data_B[4][33] ), .s(n9740), .op(
        n5815) );
  mux2_1 U12095 ( .ip1(n9814), .ip2(\cache_data_B[4][34] ), .s(n9740), .op(
        n5814) );
  mux2_1 U12096 ( .ip1(n9815), .ip2(\cache_data_B[4][35] ), .s(n9740), .op(
        n5813) );
  mux2_1 U12097 ( .ip1(n9816), .ip2(\cache_data_B[4][36] ), .s(n9740), .op(
        n5812) );
  mux2_1 U12098 ( .ip1(n9817), .ip2(\cache_data_B[4][37] ), .s(n9740), .op(
        n5811) );
  mux2_1 U12099 ( .ip1(n9818), .ip2(\cache_data_B[4][38] ), .s(n9740), .op(
        n5810) );
  mux2_1 U12100 ( .ip1(n9819), .ip2(\cache_data_B[4][39] ), .s(n9740), .op(
        n5809) );
  mux2_1 U12101 ( .ip1(n9820), .ip2(\cache_data_B[4][40] ), .s(n9740), .op(
        n5808) );
  mux2_1 U12102 ( .ip1(n9821), .ip2(\cache_data_B[4][41] ), .s(n9740), .op(
        n5807) );
  buf_1 U12103 ( .ip(n9740), .op(n9741) );
  mux2_1 U12104 ( .ip1(n9822), .ip2(\cache_data_B[4][42] ), .s(n9741), .op(
        n5806) );
  mux2_1 U12105 ( .ip1(n9823), .ip2(\cache_data_B[4][43] ), .s(n9740), .op(
        n5805) );
  mux2_1 U12106 ( .ip1(n9824), .ip2(\cache_data_B[4][44] ), .s(n9740), .op(
        n5804) );
  mux2_1 U12107 ( .ip1(n9825), .ip2(\cache_data_B[4][45] ), .s(n9740), .op(
        n5803) );
  mux2_1 U12108 ( .ip1(n9826), .ip2(\cache_data_B[4][46] ), .s(n9740), .op(
        n5802) );
  mux2_1 U12109 ( .ip1(n9827), .ip2(\cache_data_B[4][47] ), .s(n9740), .op(
        n5801) );
  mux2_1 U12110 ( .ip1(n9828), .ip2(\cache_data_B[4][48] ), .s(n9741), .op(
        n5800) );
  mux2_1 U12111 ( .ip1(n9829), .ip2(\cache_data_B[4][49] ), .s(n9741), .op(
        n5799) );
  mux2_1 U12112 ( .ip1(n9830), .ip2(\cache_data_B[4][50] ), .s(n9741), .op(
        n5798) );
  mux2_1 U12113 ( .ip1(n9831), .ip2(\cache_data_B[4][51] ), .s(n9740), .op(
        n5797) );
  mux2_1 U12114 ( .ip1(n9832), .ip2(\cache_data_B[4][52] ), .s(n9740), .op(
        n5796) );
  mux2_1 U12115 ( .ip1(n9833), .ip2(\cache_data_B[4][53] ), .s(n9740), .op(
        n5795) );
  mux2_1 U12116 ( .ip1(n9835), .ip2(\cache_data_B[4][54] ), .s(n9740), .op(
        n5794) );
  mux2_1 U12117 ( .ip1(n9836), .ip2(\cache_data_B[4][55] ), .s(n9740), .op(
        n5793) );
  mux2_1 U12118 ( .ip1(n9837), .ip2(\cache_data_B[4][56] ), .s(n9740), .op(
        n5792) );
  mux2_1 U12119 ( .ip1(n9838), .ip2(\cache_data_B[4][57] ), .s(n9741), .op(
        n5791) );
  mux2_1 U12120 ( .ip1(n9839), .ip2(\cache_data_B[4][58] ), .s(n9741), .op(
        n5790) );
  mux2_1 U12121 ( .ip1(n9840), .ip2(\cache_data_B[4][59] ), .s(n9741), .op(
        n5789) );
  mux2_1 U12122 ( .ip1(n9841), .ip2(\cache_data_B[4][60] ), .s(n9741), .op(
        n5788) );
  mux2_1 U12123 ( .ip1(n9842), .ip2(\cache_data_B[4][61] ), .s(n9741), .op(
        n5787) );
  mux2_1 U12124 ( .ip1(n9843), .ip2(\cache_data_B[4][62] ), .s(n9741), .op(
        n5786) );
  mux2_1 U12125 ( .ip1(n9845), .ip2(\cache_data_B[4][63] ), .s(n9741), .op(
        n5785) );
  nand2_1 U12126 ( .ip1(n9744), .ip2(n9807), .op(n9742) );
  mux2_1 U12127 ( .ip1(n9819), .ip2(\cache_data_B[4][71] ), .s(n9742), .op(
        n5784) );
  mux2_1 U12128 ( .ip1(n9820), .ip2(\cache_data_B[4][72] ), .s(n9742), .op(
        n5783) );
  mux2_1 U12129 ( .ip1(n9821), .ip2(\cache_data_B[4][73] ), .s(n9742), .op(
        n5782) );
  mux2_1 U12130 ( .ip1(n9822), .ip2(\cache_data_B[4][74] ), .s(n9742), .op(
        n5781) );
  mux2_1 U12131 ( .ip1(n9823), .ip2(\cache_data_B[4][75] ), .s(n9742), .op(
        n5780) );
  mux2_1 U12132 ( .ip1(n9824), .ip2(\cache_data_B[4][76] ), .s(n9742), .op(
        n5779) );
  mux2_1 U12133 ( .ip1(n9825), .ip2(\cache_data_B[4][77] ), .s(n9742), .op(
        n5778) );
  mux2_1 U12134 ( .ip1(n9826), .ip2(\cache_data_B[4][78] ), .s(n9742), .op(
        n5777) );
  buf_1 U12135 ( .ip(n9742), .op(n9743) );
  mux2_1 U12136 ( .ip1(n9827), .ip2(\cache_data_B[4][79] ), .s(n9743), .op(
        n5776) );
  mux2_1 U12137 ( .ip1(n9828), .ip2(\cache_data_B[4][80] ), .s(n9742), .op(
        n5775) );
  mux2_1 U12138 ( .ip1(n9829), .ip2(\cache_data_B[4][81] ), .s(n9742), .op(
        n5774) );
  mux2_1 U12139 ( .ip1(n9830), .ip2(\cache_data_B[4][82] ), .s(n9742), .op(
        n5773) );
  mux2_1 U12140 ( .ip1(n9831), .ip2(\cache_data_B[4][83] ), .s(n9742), .op(
        n5772) );
  mux2_1 U12141 ( .ip1(n9832), .ip2(\cache_data_B[4][84] ), .s(n9742), .op(
        n5771) );
  mux2_1 U12142 ( .ip1(n9833), .ip2(\cache_data_B[4][85] ), .s(n9742), .op(
        n5770) );
  mux2_1 U12143 ( .ip1(n9835), .ip2(\cache_data_B[4][86] ), .s(n9742), .op(
        n5769) );
  mux2_1 U12144 ( .ip1(n9836), .ip2(\cache_data_B[4][87] ), .s(n9742), .op(
        n5768) );
  mux2_1 U12145 ( .ip1(n9837), .ip2(\cache_data_B[4][88] ), .s(n9742), .op(
        n5767) );
  mux2_1 U12146 ( .ip1(n9838), .ip2(\cache_data_B[4][89] ), .s(n9743), .op(
        n5766) );
  mux2_1 U12147 ( .ip1(n9839), .ip2(\cache_data_B[4][90] ), .s(n9742), .op(
        n5765) );
  mux2_1 U12148 ( .ip1(n9840), .ip2(\cache_data_B[4][91] ), .s(n9742), .op(
        n5764) );
  mux2_1 U12149 ( .ip1(n9841), .ip2(\cache_data_B[4][92] ), .s(n9742), .op(
        n5763) );
  mux2_1 U12150 ( .ip1(n9842), .ip2(\cache_data_B[4][93] ), .s(n9742), .op(
        n5762) );
  mux2_1 U12151 ( .ip1(n9843), .ip2(\cache_data_B[4][94] ), .s(n9743), .op(
        n5761) );
  mux2_1 U12152 ( .ip1(n9845), .ip2(\cache_data_B[4][95] ), .s(n9743), .op(
        n5760) );
  mux2_1 U12153 ( .ip1(n9812), .ip2(\cache_data_B[4][64] ), .s(n9743), .op(
        n5759) );
  mux2_1 U12154 ( .ip1(n9813), .ip2(\cache_data_B[4][65] ), .s(n9743), .op(
        n5758) );
  mux2_1 U12155 ( .ip1(n9814), .ip2(\cache_data_B[4][66] ), .s(n9743), .op(
        n5757) );
  mux2_1 U12156 ( .ip1(n9815), .ip2(\cache_data_B[4][67] ), .s(n9743), .op(
        n5756) );
  mux2_1 U12157 ( .ip1(n9816), .ip2(\cache_data_B[4][68] ), .s(n9743), .op(
        n5755) );
  mux2_1 U12158 ( .ip1(n9817), .ip2(\cache_data_B[4][69] ), .s(n9743), .op(
        n5754) );
  mux2_1 U12159 ( .ip1(n9818), .ip2(\cache_data_B[4][70] ), .s(n9743), .op(
        n5753) );
  nand2_1 U12160 ( .ip1(n9744), .ip2(n9810), .op(n9745) );
  mux2_1 U12161 ( .ip1(n9812), .ip2(\cache_data_B[4][96] ), .s(n9745), .op(
        n5752) );
  mux2_1 U12162 ( .ip1(n9813), .ip2(\cache_data_B[4][97] ), .s(n9745), .op(
        n5751) );
  mux2_1 U12163 ( .ip1(n9814), .ip2(\cache_data_B[4][98] ), .s(n9745), .op(
        n5750) );
  mux2_1 U12164 ( .ip1(n9815), .ip2(\cache_data_B[4][99] ), .s(n9745), .op(
        n5749) );
  mux2_1 U12165 ( .ip1(n9816), .ip2(\cache_data_B[4][100] ), .s(n9745), .op(
        n5748) );
  mux2_1 U12166 ( .ip1(n9817), .ip2(\cache_data_B[4][101] ), .s(n9745), .op(
        n5747) );
  mux2_1 U12167 ( .ip1(n9818), .ip2(\cache_data_B[4][102] ), .s(n9745), .op(
        n5746) );
  mux2_1 U12168 ( .ip1(n9819), .ip2(\cache_data_B[4][103] ), .s(n9745), .op(
        n5745) );
  mux2_1 U12169 ( .ip1(n9820), .ip2(\cache_data_B[4][104] ), .s(n9745), .op(
        n5744) );
  mux2_1 U12170 ( .ip1(n9821), .ip2(\cache_data_B[4][105] ), .s(n9745), .op(
        n5743) );
  buf_1 U12171 ( .ip(n9745), .op(n9746) );
  mux2_1 U12172 ( .ip1(n9822), .ip2(\cache_data_B[4][106] ), .s(n9746), .op(
        n5742) );
  mux2_1 U12173 ( .ip1(n9823), .ip2(\cache_data_B[4][107] ), .s(n9745), .op(
        n5741) );
  mux2_1 U12174 ( .ip1(n9824), .ip2(\cache_data_B[4][108] ), .s(n9745), .op(
        n5740) );
  mux2_1 U12175 ( .ip1(n9825), .ip2(\cache_data_B[4][109] ), .s(n9745), .op(
        n5739) );
  mux2_1 U12176 ( .ip1(n9826), .ip2(\cache_data_B[4][110] ), .s(n9745), .op(
        n5738) );
  mux2_1 U12177 ( .ip1(n9827), .ip2(\cache_data_B[4][111] ), .s(n9745), .op(
        n5737) );
  mux2_1 U12178 ( .ip1(n9828), .ip2(\cache_data_B[4][112] ), .s(n9746), .op(
        n5736) );
  mux2_1 U12179 ( .ip1(n9829), .ip2(\cache_data_B[4][113] ), .s(n9746), .op(
        n5735) );
  mux2_1 U12180 ( .ip1(n9830), .ip2(\cache_data_B[4][114] ), .s(n9746), .op(
        n5734) );
  mux2_1 U12181 ( .ip1(n9831), .ip2(\cache_data_B[4][115] ), .s(n9745), .op(
        n5733) );
  mux2_1 U12182 ( .ip1(n9832), .ip2(\cache_data_B[4][116] ), .s(n9745), .op(
        n5732) );
  mux2_1 U12183 ( .ip1(n9833), .ip2(\cache_data_B[4][117] ), .s(n9745), .op(
        n5731) );
  mux2_1 U12184 ( .ip1(n9835), .ip2(\cache_data_B[4][118] ), .s(n9745), .op(
        n5730) );
  mux2_1 U12185 ( .ip1(n9836), .ip2(\cache_data_B[4][119] ), .s(n9745), .op(
        n5729) );
  mux2_1 U12186 ( .ip1(n9837), .ip2(\cache_data_B[4][120] ), .s(n9745), .op(
        n5728) );
  mux2_1 U12187 ( .ip1(n9838), .ip2(\cache_data_B[4][121] ), .s(n9746), .op(
        n5727) );
  mux2_1 U12188 ( .ip1(n9839), .ip2(\cache_data_B[4][122] ), .s(n9746), .op(
        n5726) );
  mux2_1 U12189 ( .ip1(n9840), .ip2(\cache_data_B[4][123] ), .s(n9746), .op(
        n5725) );
  mux2_1 U12190 ( .ip1(n9841), .ip2(\cache_data_B[4][124] ), .s(n9746), .op(
        n5724) );
  mux2_1 U12191 ( .ip1(n9842), .ip2(\cache_data_B[4][125] ), .s(n9746), .op(
        n5723) );
  mux2_1 U12192 ( .ip1(n9843), .ip2(\cache_data_B[4][126] ), .s(n9746), .op(
        n5722) );
  mux2_1 U12193 ( .ip1(n9845), .ip2(\cache_data_B[4][127] ), .s(n9746), .op(
        n5721) );
  nor2_1 U12194 ( .ip1(n9870), .ip2(n9768), .op(n9747) );
  mux2_1 U12195 ( .ip1(\cache_data_B[5][0] ), .ip2(n9770), .s(n9747), .op(
        n5720) );
  buf_1 U12196 ( .ip(n9747), .op(n9748) );
  mux2_1 U12197 ( .ip1(\cache_data_B[5][1] ), .ip2(n9813), .s(n9748), .op(
        n5719) );
  mux2_1 U12198 ( .ip1(\cache_data_B[5][2] ), .ip2(n9814), .s(n9747), .op(
        n5718) );
  mux2_1 U12199 ( .ip1(\cache_data_B[5][3] ), .ip2(n9815), .s(n9747), .op(
        n5717) );
  mux2_1 U12200 ( .ip1(\cache_data_B[5][4] ), .ip2(n9816), .s(n9747), .op(
        n5716) );
  mux2_1 U12201 ( .ip1(\cache_data_B[5][5] ), .ip2(n9817), .s(n9747), .op(
        n5715) );
  mux2_1 U12202 ( .ip1(\cache_data_B[5][6] ), .ip2(n9818), .s(n9747), .op(
        n5714) );
  mux2_1 U12203 ( .ip1(\cache_data_B[5][7] ), .ip2(n9819), .s(n9747), .op(
        n5713) );
  mux2_1 U12204 ( .ip1(\cache_data_B[5][8] ), .ip2(n9820), .s(n9747), .op(
        n5712) );
  mux2_1 U12205 ( .ip1(\cache_data_B[5][9] ), .ip2(n9821), .s(n9748), .op(
        n5711) );
  mux2_1 U12206 ( .ip1(\cache_data_B[5][10] ), .ip2(n9822), .s(n9748), .op(
        n5710) );
  mux2_1 U12207 ( .ip1(\cache_data_B[5][11] ), .ip2(n9823), .s(n9747), .op(
        n5709) );
  mux2_1 U12208 ( .ip1(\cache_data_B[5][12] ), .ip2(n9824), .s(n9747), .op(
        n5708) );
  mux2_1 U12209 ( .ip1(\cache_data_B[5][13] ), .ip2(n9825), .s(n9747), .op(
        n5707) );
  mux2_1 U12210 ( .ip1(\cache_data_B[5][14] ), .ip2(n9826), .s(n9747), .op(
        n5706) );
  mux2_1 U12211 ( .ip1(\cache_data_B[5][15] ), .ip2(n9827), .s(n9747), .op(
        n5705) );
  mux2_1 U12212 ( .ip1(\cache_data_B[5][16] ), .ip2(n9828), .s(n9747), .op(
        n5704) );
  mux2_1 U12213 ( .ip1(\cache_data_B[5][17] ), .ip2(n9787), .s(n9747), .op(
        n5703) );
  mux2_1 U12214 ( .ip1(\cache_data_B[5][18] ), .ip2(n9788), .s(n9747), .op(
        n5702) );
  mux2_1 U12215 ( .ip1(\cache_data_B[5][19] ), .ip2(n9789), .s(n9747), .op(
        n5701) );
  mux2_1 U12216 ( .ip1(\cache_data_B[5][20] ), .ip2(n9790), .s(n9747), .op(
        n5700) );
  mux2_1 U12217 ( .ip1(\cache_data_B[5][21] ), .ip2(n9791), .s(n9747), .op(
        n5699) );
  mux2_1 U12218 ( .ip1(\cache_data_B[5][22] ), .ip2(n9792), .s(n9747), .op(
        n5698) );
  mux2_1 U12219 ( .ip1(\cache_data_B[5][23] ), .ip2(n9794), .s(n9747), .op(
        n5697) );
  mux2_1 U12220 ( .ip1(\cache_data_B[5][24] ), .ip2(n9795), .s(n9748), .op(
        n5696) );
  mux2_1 U12221 ( .ip1(\cache_data_B[5][25] ), .ip2(n9796), .s(n9748), .op(
        n5695) );
  mux2_1 U12222 ( .ip1(\cache_data_B[5][26] ), .ip2(n9797), .s(n9748), .op(
        n5694) );
  mux2_1 U12223 ( .ip1(\cache_data_B[5][27] ), .ip2(n9798), .s(n9748), .op(
        n5693) );
  mux2_1 U12224 ( .ip1(\cache_data_B[5][28] ), .ip2(n9799), .s(n9748), .op(
        n5692) );
  mux2_1 U12225 ( .ip1(\cache_data_B[5][29] ), .ip2(n9800), .s(n9748), .op(
        n5691) );
  mux2_1 U12226 ( .ip1(\cache_data_B[5][30] ), .ip2(n9801), .s(n9748), .op(
        n5690) );
  mux2_1 U12227 ( .ip1(\cache_data_B[5][31] ), .ip2(n9803), .s(n9748), .op(
        n5689) );
  nand2_1 U12228 ( .ip1(n9753), .ip2(n9804), .op(n9749) );
  mux2_1 U12229 ( .ip1(n9822), .ip2(\cache_data_B[5][42] ), .s(n9749), .op(
        n5688) );
  mux2_1 U12230 ( .ip1(n9823), .ip2(\cache_data_B[5][43] ), .s(n9749), .op(
        n5687) );
  mux2_1 U12231 ( .ip1(n9824), .ip2(\cache_data_B[5][44] ), .s(n9749), .op(
        n5686) );
  mux2_1 U12232 ( .ip1(n9825), .ip2(\cache_data_B[5][45] ), .s(n9749), .op(
        n5685) );
  mux2_1 U12233 ( .ip1(n9826), .ip2(\cache_data_B[5][46] ), .s(n9749), .op(
        n5684) );
  buf_1 U12234 ( .ip(n9749), .op(n9750) );
  mux2_1 U12235 ( .ip1(n9827), .ip2(\cache_data_B[5][47] ), .s(n9750), .op(
        n5683) );
  mux2_1 U12236 ( .ip1(n9828), .ip2(\cache_data_B[5][48] ), .s(n9749), .op(
        n5682) );
  mux2_1 U12237 ( .ip1(n9829), .ip2(\cache_data_B[5][49] ), .s(n9749), .op(
        n5681) );
  mux2_1 U12238 ( .ip1(n9830), .ip2(\cache_data_B[5][50] ), .s(n9749), .op(
        n5680) );
  mux2_1 U12239 ( .ip1(n9831), .ip2(\cache_data_B[5][51] ), .s(n9749), .op(
        n5679) );
  mux2_1 U12240 ( .ip1(n9832), .ip2(\cache_data_B[5][52] ), .s(n9749), .op(
        n5678) );
  mux2_1 U12241 ( .ip1(n9833), .ip2(\cache_data_B[5][53] ), .s(n9749), .op(
        n5677) );
  mux2_1 U12242 ( .ip1(n9835), .ip2(\cache_data_B[5][54] ), .s(n9749), .op(
        n5676) );
  mux2_1 U12243 ( .ip1(n9836), .ip2(\cache_data_B[5][55] ), .s(n9749), .op(
        n5675) );
  mux2_1 U12244 ( .ip1(n9837), .ip2(\cache_data_B[5][56] ), .s(n9749), .op(
        n5674) );
  mux2_1 U12245 ( .ip1(n9838), .ip2(\cache_data_B[5][57] ), .s(n9750), .op(
        n5673) );
  mux2_1 U12246 ( .ip1(n9839), .ip2(\cache_data_B[5][58] ), .s(n9749), .op(
        n5672) );
  mux2_1 U12247 ( .ip1(n9840), .ip2(\cache_data_B[5][59] ), .s(n9749), .op(
        n5671) );
  mux2_1 U12248 ( .ip1(n9841), .ip2(\cache_data_B[5][60] ), .s(n9749), .op(
        n5670) );
  mux2_1 U12249 ( .ip1(n9842), .ip2(\cache_data_B[5][61] ), .s(n9749), .op(
        n5669) );
  mux2_1 U12250 ( .ip1(n9843), .ip2(\cache_data_B[5][62] ), .s(n9749), .op(
        n5668) );
  mux2_1 U12251 ( .ip1(n9845), .ip2(\cache_data_B[5][63] ), .s(n9749), .op(
        n5667) );
  mux2_1 U12252 ( .ip1(n9812), .ip2(\cache_data_B[5][32] ), .s(n9749), .op(
        n5666) );
  mux2_1 U12253 ( .ip1(n9813), .ip2(\cache_data_B[5][33] ), .s(n9750), .op(
        n5665) );
  mux2_1 U12254 ( .ip1(n9814), .ip2(\cache_data_B[5][34] ), .s(n9750), .op(
        n5664) );
  mux2_1 U12255 ( .ip1(n9815), .ip2(\cache_data_B[5][35] ), .s(n9750), .op(
        n5663) );
  mux2_1 U12256 ( .ip1(n9816), .ip2(\cache_data_B[5][36] ), .s(n9750), .op(
        n5662) );
  mux2_1 U12257 ( .ip1(n9817), .ip2(\cache_data_B[5][37] ), .s(n9750), .op(
        n5661) );
  mux2_1 U12258 ( .ip1(n9818), .ip2(\cache_data_B[5][38] ), .s(n9750), .op(
        n5660) );
  mux2_1 U12259 ( .ip1(n9819), .ip2(\cache_data_B[5][39] ), .s(n9750), .op(
        n5659) );
  mux2_1 U12260 ( .ip1(n9820), .ip2(\cache_data_B[5][40] ), .s(n9750), .op(
        n5658) );
  mux2_1 U12261 ( .ip1(n9821), .ip2(\cache_data_B[5][41] ), .s(n9750), .op(
        n5657) );
  nor2_1 U12262 ( .ip1(n9870), .ip2(n9761), .op(n9751) );
  buf_1 U12263 ( .ip(n9751), .op(n9752) );
  mux2_1 U12264 ( .ip1(\cache_data_B[5][64] ), .ip2(n9812), .s(n9752), .op(
        n5656) );
  mux2_1 U12265 ( .ip1(\cache_data_B[5][65] ), .ip2(n9771), .s(n9751), .op(
        n5655) );
  mux2_1 U12266 ( .ip1(\cache_data_B[5][66] ), .ip2(n9772), .s(n9751), .op(
        n5654) );
  mux2_1 U12267 ( .ip1(\cache_data_B[5][67] ), .ip2(n9773), .s(n9751), .op(
        n5653) );
  mux2_1 U12268 ( .ip1(\cache_data_B[5][68] ), .ip2(n9774), .s(n9751), .op(
        n5652) );
  mux2_1 U12269 ( .ip1(\cache_data_B[5][69] ), .ip2(n9775), .s(n9751), .op(
        n5651) );
  mux2_1 U12270 ( .ip1(\cache_data_B[5][70] ), .ip2(n9776), .s(n9751), .op(
        n5650) );
  mux2_1 U12271 ( .ip1(\cache_data_B[5][71] ), .ip2(n9777), .s(n9751), .op(
        n5649) );
  mux2_1 U12272 ( .ip1(\cache_data_B[5][72] ), .ip2(n9778), .s(n9751), .op(
        n5648) );
  mux2_1 U12273 ( .ip1(\cache_data_B[5][73] ), .ip2(n9779), .s(n9752), .op(
        n5647) );
  mux2_1 U12274 ( .ip1(\cache_data_B[5][74] ), .ip2(n9780), .s(n9752), .op(
        n5646) );
  mux2_1 U12275 ( .ip1(\cache_data_B[5][75] ), .ip2(n9781), .s(n9751), .op(
        n5645) );
  mux2_1 U12276 ( .ip1(\cache_data_B[5][76] ), .ip2(n9782), .s(n9751), .op(
        n5644) );
  mux2_1 U12277 ( .ip1(\cache_data_B[5][77] ), .ip2(n9783), .s(n9751), .op(
        n5643) );
  mux2_1 U12278 ( .ip1(\cache_data_B[5][78] ), .ip2(n9784), .s(n9751), .op(
        n5642) );
  mux2_1 U12279 ( .ip1(\cache_data_B[5][79] ), .ip2(n9785), .s(n9751), .op(
        n5641) );
  mux2_1 U12280 ( .ip1(\cache_data_B[5][80] ), .ip2(n9786), .s(n9751), .op(
        n5640) );
  mux2_1 U12281 ( .ip1(\cache_data_B[5][81] ), .ip2(n9829), .s(n9751), .op(
        n5639) );
  mux2_1 U12282 ( .ip1(\cache_data_B[5][82] ), .ip2(n9830), .s(n9751), .op(
        n5638) );
  mux2_1 U12283 ( .ip1(\cache_data_B[5][83] ), .ip2(n9789), .s(n9751), .op(
        n5637) );
  mux2_1 U12284 ( .ip1(\cache_data_B[5][84] ), .ip2(n9790), .s(n9751), .op(
        n5636) );
  mux2_1 U12285 ( .ip1(\cache_data_B[5][85] ), .ip2(n9791), .s(n9751), .op(
        n5635) );
  mux2_1 U12286 ( .ip1(\cache_data_B[5][86] ), .ip2(n9792), .s(n9751), .op(
        n5634) );
  mux2_1 U12287 ( .ip1(\cache_data_B[5][87] ), .ip2(n9794), .s(n9751), .op(
        n5633) );
  mux2_1 U12288 ( .ip1(\cache_data_B[5][88] ), .ip2(n9795), .s(n9752), .op(
        n5632) );
  mux2_1 U12289 ( .ip1(\cache_data_B[5][89] ), .ip2(n9838), .s(n9752), .op(
        n5631) );
  mux2_1 U12290 ( .ip1(\cache_data_B[5][90] ), .ip2(n9839), .s(n9752), .op(
        n5630) );
  mux2_1 U12291 ( .ip1(\cache_data_B[5][91] ), .ip2(n9840), .s(n9752), .op(
        n5629) );
  mux2_1 U12292 ( .ip1(\cache_data_B[5][92] ), .ip2(n9841), .s(n9752), .op(
        n5628) );
  mux2_1 U12293 ( .ip1(\cache_data_B[5][93] ), .ip2(n9842), .s(n9752), .op(
        n5627) );
  mux2_1 U12294 ( .ip1(\cache_data_B[5][94] ), .ip2(n9843), .s(n9752), .op(
        n5626) );
  mux2_1 U12295 ( .ip1(\cache_data_B[5][95] ), .ip2(n9845), .s(n9752), .op(
        n5625) );
  nand2_1 U12296 ( .ip1(n9753), .ip2(n9810), .op(n9754) );
  mux2_1 U12297 ( .ip1(n9812), .ip2(\cache_data_B[5][96] ), .s(n9754), .op(
        n5624) );
  mux2_1 U12298 ( .ip1(n9813), .ip2(\cache_data_B[5][97] ), .s(n9754), .op(
        n5623) );
  mux2_1 U12299 ( .ip1(n9814), .ip2(\cache_data_B[5][98] ), .s(n9754), .op(
        n5622) );
  mux2_1 U12300 ( .ip1(n9815), .ip2(\cache_data_B[5][99] ), .s(n9754), .op(
        n5621) );
  mux2_1 U12301 ( .ip1(n9816), .ip2(\cache_data_B[5][100] ), .s(n9754), .op(
        n5620) );
  mux2_1 U12302 ( .ip1(n9817), .ip2(\cache_data_B[5][101] ), .s(n9754), .op(
        n5619) );
  mux2_1 U12303 ( .ip1(n9818), .ip2(\cache_data_B[5][102] ), .s(n9754), .op(
        n5618) );
  mux2_1 U12304 ( .ip1(n9819), .ip2(\cache_data_B[5][103] ), .s(n9754), .op(
        n5617) );
  mux2_1 U12305 ( .ip1(n9820), .ip2(\cache_data_B[5][104] ), .s(n9754), .op(
        n5616) );
  mux2_1 U12306 ( .ip1(n9821), .ip2(\cache_data_B[5][105] ), .s(n9754), .op(
        n5615) );
  buf_1 U12307 ( .ip(n9754), .op(n9755) );
  mux2_1 U12308 ( .ip1(n9822), .ip2(\cache_data_B[5][106] ), .s(n9755), .op(
        n5614) );
  mux2_1 U12309 ( .ip1(n9823), .ip2(\cache_data_B[5][107] ), .s(n9754), .op(
        n5613) );
  mux2_1 U12310 ( .ip1(n9824), .ip2(\cache_data_B[5][108] ), .s(n9754), .op(
        n5612) );
  mux2_1 U12311 ( .ip1(n9825), .ip2(\cache_data_B[5][109] ), .s(n9754), .op(
        n5611) );
  mux2_1 U12312 ( .ip1(n9826), .ip2(\cache_data_B[5][110] ), .s(n9754), .op(
        n5610) );
  mux2_1 U12313 ( .ip1(n9827), .ip2(\cache_data_B[5][111] ), .s(n9754), .op(
        n5609) );
  mux2_1 U12314 ( .ip1(n9828), .ip2(\cache_data_B[5][112] ), .s(n9755), .op(
        n5608) );
  mux2_1 U12315 ( .ip1(n9829), .ip2(\cache_data_B[5][113] ), .s(n9755), .op(
        n5607) );
  mux2_1 U12316 ( .ip1(n9830), .ip2(\cache_data_B[5][114] ), .s(n9755), .op(
        n5606) );
  mux2_1 U12317 ( .ip1(n9831), .ip2(\cache_data_B[5][115] ), .s(n9754), .op(
        n5605) );
  mux2_1 U12318 ( .ip1(n9832), .ip2(\cache_data_B[5][116] ), .s(n9754), .op(
        n5604) );
  mux2_1 U12319 ( .ip1(n9833), .ip2(\cache_data_B[5][117] ), .s(n9754), .op(
        n5603) );
  mux2_1 U12320 ( .ip1(n9835), .ip2(\cache_data_B[5][118] ), .s(n9754), .op(
        n5602) );
  mux2_1 U12321 ( .ip1(n9836), .ip2(\cache_data_B[5][119] ), .s(n9754), .op(
        n5601) );
  mux2_1 U12322 ( .ip1(n9837), .ip2(\cache_data_B[5][120] ), .s(n9754), .op(
        n5600) );
  mux2_1 U12323 ( .ip1(n9838), .ip2(\cache_data_B[5][121] ), .s(n9755), .op(
        n5599) );
  mux2_1 U12324 ( .ip1(n9839), .ip2(\cache_data_B[5][122] ), .s(n9755), .op(
        n5598) );
  mux2_1 U12325 ( .ip1(n9840), .ip2(\cache_data_B[5][123] ), .s(n9755), .op(
        n5597) );
  mux2_1 U12326 ( .ip1(n9841), .ip2(\cache_data_B[5][124] ), .s(n9755), .op(
        n5596) );
  mux2_1 U12327 ( .ip1(n9842), .ip2(\cache_data_B[5][125] ), .s(n9755), .op(
        n5595) );
  mux2_1 U12328 ( .ip1(n9843), .ip2(\cache_data_B[5][126] ), .s(n9755), .op(
        n5594) );
  mux2_1 U12329 ( .ip1(n9845), .ip2(\cache_data_B[5][127] ), .s(n9755), .op(
        n5593) );
  nand2_1 U12330 ( .ip1(n9765), .ip2(n9756), .op(n9757) );
  mux2_1 U12331 ( .ip1(n9825), .ip2(\cache_data_B[6][13] ), .s(n9757), .op(
        n5592) );
  mux2_1 U12332 ( .ip1(n9826), .ip2(\cache_data_B[6][14] ), .s(n9757), .op(
        n5591) );
  mux2_1 U12333 ( .ip1(n9827), .ip2(\cache_data_B[6][15] ), .s(n9757), .op(
        n5590) );
  mux2_1 U12334 ( .ip1(n9828), .ip2(\cache_data_B[6][16] ), .s(n9757), .op(
        n5589) );
  mux2_1 U12335 ( .ip1(n9829), .ip2(\cache_data_B[6][17] ), .s(n9757), .op(
        n5588) );
  mux2_1 U12336 ( .ip1(n9830), .ip2(\cache_data_B[6][18] ), .s(n9757), .op(
        n5587) );
  mux2_1 U12337 ( .ip1(n9831), .ip2(\cache_data_B[6][19] ), .s(n9757), .op(
        n5586) );
  mux2_1 U12338 ( .ip1(n9832), .ip2(\cache_data_B[6][20] ), .s(n9757), .op(
        n5585) );
  mux2_1 U12339 ( .ip1(n9833), .ip2(\cache_data_B[6][21] ), .s(n9757), .op(
        n5584) );
  mux2_1 U12340 ( .ip1(n9835), .ip2(\cache_data_B[6][22] ), .s(n9757), .op(
        n5583) );
  mux2_1 U12341 ( .ip1(n9836), .ip2(\cache_data_B[6][23] ), .s(n9757), .op(
        n5582) );
  mux2_1 U12342 ( .ip1(n9837), .ip2(\cache_data_B[6][24] ), .s(n9757), .op(
        n5581) );
  mux2_1 U12343 ( .ip1(n9838), .ip2(\cache_data_B[6][25] ), .s(n9757), .op(
        n5580) );
  mux2_1 U12344 ( .ip1(n9839), .ip2(\cache_data_B[6][26] ), .s(n9757), .op(
        n5579) );
  mux2_1 U12345 ( .ip1(n9840), .ip2(\cache_data_B[6][27] ), .s(n9757), .op(
        n5578) );
  mux2_1 U12346 ( .ip1(n9841), .ip2(\cache_data_B[6][28] ), .s(n9757), .op(
        n5577) );
  mux2_1 U12347 ( .ip1(n9842), .ip2(\cache_data_B[6][29] ), .s(n9757), .op(
        n5576) );
  mux2_1 U12348 ( .ip1(n9843), .ip2(\cache_data_B[6][30] ), .s(n9757), .op(
        n5575) );
  buf_1 U12349 ( .ip(n9757), .op(n9758) );
  mux2_1 U12350 ( .ip1(n9845), .ip2(\cache_data_B[6][31] ), .s(n9758), .op(
        n5574) );
  mux2_1 U12351 ( .ip1(n9812), .ip2(\cache_data_B[6][0] ), .s(n9758), .op(
        n5573) );
  mux2_1 U12352 ( .ip1(n9813), .ip2(\cache_data_B[6][1] ), .s(n9758), .op(
        n5572) );
  mux2_1 U12353 ( .ip1(n9814), .ip2(\cache_data_B[6][2] ), .s(n9758), .op(
        n5571) );
  mux2_1 U12354 ( .ip1(n9815), .ip2(\cache_data_B[6][3] ), .s(n9758), .op(
        n5570) );
  mux2_1 U12355 ( .ip1(n9816), .ip2(\cache_data_B[6][4] ), .s(n9757), .op(
        n5569) );
  mux2_1 U12356 ( .ip1(n9817), .ip2(\cache_data_B[6][5] ), .s(n9757), .op(
        n5568) );
  mux2_1 U12357 ( .ip1(n9818), .ip2(\cache_data_B[6][6] ), .s(n9757), .op(
        n5567) );
  mux2_1 U12358 ( .ip1(n9819), .ip2(\cache_data_B[6][7] ), .s(n9758), .op(
        n5566) );
  mux2_1 U12359 ( .ip1(n9820), .ip2(\cache_data_B[6][8] ), .s(n9758), .op(
        n5565) );
  mux2_1 U12360 ( .ip1(n9821), .ip2(\cache_data_B[6][9] ), .s(n9758), .op(
        n5564) );
  mux2_1 U12361 ( .ip1(n9822), .ip2(\cache_data_B[6][10] ), .s(n9758), .op(
        n5563) );
  mux2_1 U12362 ( .ip1(n9823), .ip2(\cache_data_B[6][11] ), .s(n9758), .op(
        n5562) );
  mux2_1 U12363 ( .ip1(n9824), .ip2(\cache_data_B[6][12] ), .s(n9758), .op(
        n5561) );
  nand2_1 U12364 ( .ip1(n9765), .ip2(n9804), .op(n9759) );
  mux2_1 U12365 ( .ip1(n9812), .ip2(\cache_data_B[6][32] ), .s(n9759), .op(
        n5560) );
  mux2_1 U12366 ( .ip1(n9813), .ip2(\cache_data_B[6][33] ), .s(n9759), .op(
        n5559) );
  mux2_1 U12367 ( .ip1(n9814), .ip2(\cache_data_B[6][34] ), .s(n9759), .op(
        n5558) );
  mux2_1 U12368 ( .ip1(n9815), .ip2(\cache_data_B[6][35] ), .s(n9759), .op(
        n5557) );
  mux2_1 U12369 ( .ip1(n9816), .ip2(\cache_data_B[6][36] ), .s(n9759), .op(
        n5556) );
  mux2_1 U12370 ( .ip1(n9817), .ip2(\cache_data_B[6][37] ), .s(n9759), .op(
        n5555) );
  mux2_1 U12371 ( .ip1(n9818), .ip2(\cache_data_B[6][38] ), .s(n9759), .op(
        n5554) );
  mux2_1 U12372 ( .ip1(n9819), .ip2(\cache_data_B[6][39] ), .s(n9759), .op(
        n5553) );
  mux2_1 U12373 ( .ip1(n9820), .ip2(\cache_data_B[6][40] ), .s(n9759), .op(
        n5552) );
  mux2_1 U12374 ( .ip1(n9821), .ip2(\cache_data_B[6][41] ), .s(n9759), .op(
        n5551) );
  buf_1 U12375 ( .ip(n9759), .op(n9760) );
  mux2_1 U12376 ( .ip1(n9822), .ip2(\cache_data_B[6][42] ), .s(n9760), .op(
        n5550) );
  mux2_1 U12377 ( .ip1(n9823), .ip2(\cache_data_B[6][43] ), .s(n9759), .op(
        n5549) );
  mux2_1 U12378 ( .ip1(n9824), .ip2(\cache_data_B[6][44] ), .s(n9759), .op(
        n5548) );
  mux2_1 U12379 ( .ip1(n9825), .ip2(\cache_data_B[6][45] ), .s(n9759), .op(
        n5547) );
  mux2_1 U12380 ( .ip1(n9826), .ip2(\cache_data_B[6][46] ), .s(n9759), .op(
        n5546) );
  mux2_1 U12381 ( .ip1(n9827), .ip2(\cache_data_B[6][47] ), .s(n9759), .op(
        n5545) );
  mux2_1 U12382 ( .ip1(n9828), .ip2(\cache_data_B[6][48] ), .s(n9760), .op(
        n5544) );
  mux2_1 U12383 ( .ip1(n9829), .ip2(\cache_data_B[6][49] ), .s(n9760), .op(
        n5543) );
  mux2_1 U12384 ( .ip1(n9830), .ip2(\cache_data_B[6][50] ), .s(n9760), .op(
        n5542) );
  mux2_1 U12385 ( .ip1(n9831), .ip2(\cache_data_B[6][51] ), .s(n9759), .op(
        n5541) );
  mux2_1 U12386 ( .ip1(n9832), .ip2(\cache_data_B[6][52] ), .s(n9759), .op(
        n5540) );
  mux2_1 U12387 ( .ip1(n9833), .ip2(\cache_data_B[6][53] ), .s(n9759), .op(
        n5539) );
  mux2_1 U12388 ( .ip1(n9835), .ip2(\cache_data_B[6][54] ), .s(n9759), .op(
        n5538) );
  mux2_1 U12389 ( .ip1(n9836), .ip2(\cache_data_B[6][55] ), .s(n9759), .op(
        n5537) );
  mux2_1 U12390 ( .ip1(n9837), .ip2(\cache_data_B[6][56] ), .s(n9759), .op(
        n5536) );
  mux2_1 U12391 ( .ip1(n9838), .ip2(\cache_data_B[6][57] ), .s(n9760), .op(
        n5535) );
  mux2_1 U12392 ( .ip1(n9839), .ip2(\cache_data_B[6][58] ), .s(n9760), .op(
        n5534) );
  mux2_1 U12393 ( .ip1(n9840), .ip2(\cache_data_B[6][59] ), .s(n9760), .op(
        n5533) );
  mux2_1 U12394 ( .ip1(n9841), .ip2(\cache_data_B[6][60] ), .s(n9760), .op(
        n5532) );
  mux2_1 U12395 ( .ip1(n9842), .ip2(\cache_data_B[6][61] ), .s(n9760), .op(
        n5531) );
  mux2_1 U12396 ( .ip1(n9843), .ip2(\cache_data_B[6][62] ), .s(n9760), .op(
        n5530) );
  mux2_1 U12397 ( .ip1(n9845), .ip2(\cache_data_B[6][63] ), .s(n9760), .op(
        n5529) );
  nor2_1 U12398 ( .ip1(n9762), .ip2(n9761), .op(n9763) );
  buf_1 U12399 ( .ip(n9763), .op(n9764) );
  mux2_1 U12400 ( .ip1(\cache_data_B[6][64] ), .ip2(n9770), .s(n9764), .op(
        n5528) );
  mux2_1 U12401 ( .ip1(\cache_data_B[6][65] ), .ip2(n9771), .s(n9763), .op(
        n5527) );
  mux2_1 U12402 ( .ip1(\cache_data_B[6][66] ), .ip2(n9772), .s(n9763), .op(
        n5526) );
  mux2_1 U12403 ( .ip1(\cache_data_B[6][67] ), .ip2(n9773), .s(n9763), .op(
        n5525) );
  mux2_1 U12404 ( .ip1(\cache_data_B[6][68] ), .ip2(n9774), .s(n9763), .op(
        n5524) );
  mux2_1 U12405 ( .ip1(\cache_data_B[6][69] ), .ip2(n9775), .s(n9763), .op(
        n5523) );
  mux2_1 U12406 ( .ip1(\cache_data_B[6][70] ), .ip2(n9776), .s(n9763), .op(
        n5522) );
  mux2_1 U12407 ( .ip1(\cache_data_B[6][71] ), .ip2(n9777), .s(n9763), .op(
        n5521) );
  mux2_1 U12408 ( .ip1(\cache_data_B[6][72] ), .ip2(n9778), .s(n9763), .op(
        n5520) );
  mux2_1 U12409 ( .ip1(\cache_data_B[6][73] ), .ip2(n9779), .s(n9763), .op(
        n5519) );
  mux2_1 U12410 ( .ip1(\cache_data_B[6][74] ), .ip2(n9780), .s(n9763), .op(
        n5518) );
  mux2_1 U12411 ( .ip1(\cache_data_B[6][75] ), .ip2(n9781), .s(n9763), .op(
        n5517) );
  mux2_1 U12412 ( .ip1(\cache_data_B[6][76] ), .ip2(n9782), .s(n9763), .op(
        n5516) );
  mux2_1 U12413 ( .ip1(\cache_data_B[6][77] ), .ip2(n9783), .s(n9763), .op(
        n5515) );
  mux2_1 U12414 ( .ip1(\cache_data_B[6][78] ), .ip2(n9784), .s(n9763), .op(
        n5514) );
  mux2_1 U12415 ( .ip1(\cache_data_B[6][79] ), .ip2(n9785), .s(n9763), .op(
        n5513) );
  mux2_1 U12416 ( .ip1(\cache_data_B[6][80] ), .ip2(n9786), .s(n9763), .op(
        n5512) );
  mux2_1 U12417 ( .ip1(\cache_data_B[6][81] ), .ip2(n9787), .s(n9763), .op(
        n5511) );
  mux2_1 U12418 ( .ip1(\cache_data_B[6][82] ), .ip2(n9788), .s(n9763), .op(
        n5510) );
  mux2_1 U12419 ( .ip1(\cache_data_B[6][83] ), .ip2(n9789), .s(n9763), .op(
        n5509) );
  mux2_1 U12420 ( .ip1(\cache_data_B[6][84] ), .ip2(n9790), .s(n9764), .op(
        n5508) );
  mux2_1 U12421 ( .ip1(\cache_data_B[6][85] ), .ip2(n9791), .s(n9764), .op(
        n5507) );
  mux2_1 U12422 ( .ip1(\cache_data_B[6][86] ), .ip2(n9792), .s(n9764), .op(
        n5506) );
  mux2_1 U12423 ( .ip1(\cache_data_B[6][87] ), .ip2(n9794), .s(n9764), .op(
        n5505) );
  mux2_1 U12424 ( .ip1(\cache_data_B[6][88] ), .ip2(n9795), .s(n9763), .op(
        n5504) );
  mux2_1 U12425 ( .ip1(\cache_data_B[6][89] ), .ip2(n9796), .s(n9763), .op(
        n5503) );
  mux2_1 U12426 ( .ip1(\cache_data_B[6][90] ), .ip2(n9797), .s(n9764), .op(
        n5502) );
  mux2_1 U12427 ( .ip1(\cache_data_B[6][91] ), .ip2(n9798), .s(n9764), .op(
        n5501) );
  mux2_1 U12428 ( .ip1(\cache_data_B[6][92] ), .ip2(n9799), .s(n9764), .op(
        n5500) );
  mux2_1 U12429 ( .ip1(\cache_data_B[6][93] ), .ip2(n9800), .s(n9764), .op(
        n5499) );
  mux2_1 U12430 ( .ip1(\cache_data_B[6][94] ), .ip2(n9801), .s(n9764), .op(
        n5498) );
  mux2_1 U12431 ( .ip1(\cache_data_B[6][95] ), .ip2(n9803), .s(n9764), .op(
        n5497) );
  nand2_1 U12432 ( .ip1(n9765), .ip2(n9810), .op(n9766) );
  mux2_1 U12433 ( .ip1(n9828), .ip2(\cache_data_B[6][112] ), .s(n9766), .op(
        n5496) );
  mux2_1 U12434 ( .ip1(n9829), .ip2(\cache_data_B[6][113] ), .s(n9766), .op(
        n5495) );
  mux2_1 U12435 ( .ip1(n9830), .ip2(\cache_data_B[6][114] ), .s(n9766), .op(
        n5494) );
  mux2_1 U12436 ( .ip1(n9831), .ip2(\cache_data_B[6][115] ), .s(n9766), .op(
        n5493) );
  mux2_1 U12437 ( .ip1(n9832), .ip2(\cache_data_B[6][116] ), .s(n9766), .op(
        n5492) );
  mux2_1 U12438 ( .ip1(n9833), .ip2(\cache_data_B[6][117] ), .s(n9766), .op(
        n5491) );
  mux2_1 U12439 ( .ip1(n9835), .ip2(\cache_data_B[6][118] ), .s(n9766), .op(
        n5490) );
  mux2_1 U12440 ( .ip1(n9836), .ip2(\cache_data_B[6][119] ), .s(n9766), .op(
        n5489) );
  mux2_1 U12441 ( .ip1(n9837), .ip2(\cache_data_B[6][120] ), .s(n9766), .op(
        n5488) );
  mux2_1 U12442 ( .ip1(n9838), .ip2(\cache_data_B[6][121] ), .s(n9766), .op(
        n5487) );
  mux2_1 U12443 ( .ip1(n9839), .ip2(\cache_data_B[6][122] ), .s(n9766), .op(
        n5486) );
  mux2_1 U12444 ( .ip1(n9840), .ip2(\cache_data_B[6][123] ), .s(n9766), .op(
        n5485) );
  mux2_1 U12445 ( .ip1(n9841), .ip2(\cache_data_B[6][124] ), .s(n9766), .op(
        n5484) );
  mux2_1 U12446 ( .ip1(n9842), .ip2(\cache_data_B[6][125] ), .s(n9766), .op(
        n5483) );
  mux2_1 U12447 ( .ip1(n9843), .ip2(\cache_data_B[6][126] ), .s(n9766), .op(
        n5482) );
  mux2_1 U12448 ( .ip1(n9845), .ip2(\cache_data_B[6][127] ), .s(n9766), .op(
        n5481) );
  mux2_1 U12449 ( .ip1(n9812), .ip2(\cache_data_B[6][96] ), .s(n9766), .op(
        n5480) );
  mux2_1 U12450 ( .ip1(n9813), .ip2(\cache_data_B[6][97] ), .s(n9766), .op(
        n5479) );
  buf_1 U12451 ( .ip(n9766), .op(n9767) );
  mux2_1 U12452 ( .ip1(n9814), .ip2(\cache_data_B[6][98] ), .s(n9767), .op(
        n5478) );
  mux2_1 U12453 ( .ip1(n9815), .ip2(\cache_data_B[6][99] ), .s(n9767), .op(
        n5477) );
  mux2_1 U12454 ( .ip1(n9816), .ip2(\cache_data_B[6][100] ), .s(n9766), .op(
        n5476) );
  mux2_1 U12455 ( .ip1(n9817), .ip2(\cache_data_B[6][101] ), .s(n9767), .op(
        n5475) );
  mux2_1 U12456 ( .ip1(n9818), .ip2(\cache_data_B[6][102] ), .s(n9767), .op(
        n5474) );
  mux2_1 U12457 ( .ip1(n9819), .ip2(\cache_data_B[6][103] ), .s(n9767), .op(
        n5473) );
  mux2_1 U12458 ( .ip1(n9820), .ip2(\cache_data_B[6][104] ), .s(n9766), .op(
        n5472) );
  mux2_1 U12459 ( .ip1(n9821), .ip2(\cache_data_B[6][105] ), .s(n9766), .op(
        n5471) );
  mux2_1 U12460 ( .ip1(n9822), .ip2(\cache_data_B[6][106] ), .s(n9767), .op(
        n5470) );
  mux2_1 U12461 ( .ip1(n9823), .ip2(\cache_data_B[6][107] ), .s(n9767), .op(
        n5469) );
  mux2_1 U12462 ( .ip1(n9824), .ip2(\cache_data_B[6][108] ), .s(n9767), .op(
        n5468) );
  mux2_1 U12463 ( .ip1(n9825), .ip2(\cache_data_B[6][109] ), .s(n9767), .op(
        n5467) );
  mux2_1 U12464 ( .ip1(n9826), .ip2(\cache_data_B[6][110] ), .s(n9767), .op(
        n5466) );
  mux2_1 U12465 ( .ip1(n9827), .ip2(\cache_data_B[6][111] ), .s(n9767), .op(
        n5465) );
  nor2_1 U12466 ( .ip1(n9769), .ip2(n9768), .op(n9793) );
  buf_1 U12467 ( .ip(n9793), .op(n9802) );
  mux2_1 U12468 ( .ip1(\cache_data_B[7][0] ), .ip2(n9770), .s(n9802), .op(
        n5464) );
  mux2_1 U12469 ( .ip1(\cache_data_B[7][1] ), .ip2(n9771), .s(n9793), .op(
        n5463) );
  mux2_1 U12470 ( .ip1(\cache_data_B[7][2] ), .ip2(n9772), .s(n9793), .op(
        n5462) );
  mux2_1 U12471 ( .ip1(\cache_data_B[7][3] ), .ip2(n9773), .s(n9793), .op(
        n5461) );
  mux2_1 U12472 ( .ip1(\cache_data_B[7][4] ), .ip2(n9774), .s(n9793), .op(
        n5460) );
  mux2_1 U12473 ( .ip1(\cache_data_B[7][5] ), .ip2(n9775), .s(n9793), .op(
        n5459) );
  mux2_1 U12474 ( .ip1(\cache_data_B[7][6] ), .ip2(n9776), .s(n9793), .op(
        n5458) );
  mux2_1 U12475 ( .ip1(\cache_data_B[7][7] ), .ip2(n9777), .s(n9793), .op(
        n5457) );
  mux2_1 U12476 ( .ip1(\cache_data_B[7][8] ), .ip2(n9778), .s(n9793), .op(
        n5456) );
  mux2_1 U12477 ( .ip1(\cache_data_B[7][9] ), .ip2(n9779), .s(n9802), .op(
        n5455) );
  mux2_1 U12478 ( .ip1(\cache_data_B[7][10] ), .ip2(n9780), .s(n9802), .op(
        n5454) );
  mux2_1 U12479 ( .ip1(\cache_data_B[7][11] ), .ip2(n9781), .s(n9793), .op(
        n5453) );
  mux2_1 U12480 ( .ip1(\cache_data_B[7][12] ), .ip2(n9782), .s(n9793), .op(
        n5452) );
  mux2_1 U12481 ( .ip1(\cache_data_B[7][13] ), .ip2(n9783), .s(n9793), .op(
        n5451) );
  mux2_1 U12482 ( .ip1(\cache_data_B[7][14] ), .ip2(n9784), .s(n9793), .op(
        n5450) );
  mux2_1 U12483 ( .ip1(\cache_data_B[7][15] ), .ip2(n9785), .s(n9793), .op(
        n5449) );
  mux2_1 U12484 ( .ip1(\cache_data_B[7][16] ), .ip2(n9786), .s(n9793), .op(
        n5448) );
  mux2_1 U12485 ( .ip1(\cache_data_B[7][17] ), .ip2(n9787), .s(n9793), .op(
        n5447) );
  mux2_1 U12486 ( .ip1(\cache_data_B[7][18] ), .ip2(n9788), .s(n9793), .op(
        n5446) );
  mux2_1 U12487 ( .ip1(\cache_data_B[7][19] ), .ip2(n9789), .s(n9793), .op(
        n5445) );
  mux2_1 U12488 ( .ip1(\cache_data_B[7][20] ), .ip2(n9790), .s(n9793), .op(
        n5444) );
  mux2_1 U12489 ( .ip1(\cache_data_B[7][21] ), .ip2(n9791), .s(n9793), .op(
        n5443) );
  mux2_1 U12490 ( .ip1(\cache_data_B[7][22] ), .ip2(n9792), .s(n9793), .op(
        n5442) );
  mux2_1 U12491 ( .ip1(\cache_data_B[7][23] ), .ip2(n9794), .s(n9793), .op(
        n5441) );
  mux2_1 U12492 ( .ip1(\cache_data_B[7][24] ), .ip2(n9795), .s(n9802), .op(
        n5440) );
  mux2_1 U12493 ( .ip1(\cache_data_B[7][25] ), .ip2(n9796), .s(n9802), .op(
        n5439) );
  mux2_1 U12494 ( .ip1(\cache_data_B[7][26] ), .ip2(n9797), .s(n9802), .op(
        n5438) );
  mux2_1 U12495 ( .ip1(\cache_data_B[7][27] ), .ip2(n9798), .s(n9802), .op(
        n5437) );
  mux2_1 U12496 ( .ip1(\cache_data_B[7][28] ), .ip2(n9799), .s(n9802), .op(
        n5436) );
  mux2_1 U12497 ( .ip1(\cache_data_B[7][29] ), .ip2(n9800), .s(n9802), .op(
        n5435) );
  mux2_1 U12498 ( .ip1(\cache_data_B[7][30] ), .ip2(n9801), .s(n9802), .op(
        n5434) );
  mux2_1 U12499 ( .ip1(\cache_data_B[7][31] ), .ip2(n9803), .s(n9802), .op(
        n5433) );
  nand2_1 U12500 ( .ip1(n9811), .ip2(n9804), .op(n9805) );
  mux2_1 U12501 ( .ip1(n9812), .ip2(\cache_data_B[7][32] ), .s(n9805), .op(
        n5432) );
  mux2_1 U12502 ( .ip1(n9813), .ip2(\cache_data_B[7][33] ), .s(n9805), .op(
        n5431) );
  mux2_1 U12503 ( .ip1(n9814), .ip2(\cache_data_B[7][34] ), .s(n9805), .op(
        n5430) );
  mux2_1 U12504 ( .ip1(n9815), .ip2(\cache_data_B[7][35] ), .s(n9805), .op(
        n5429) );
  mux2_1 U12505 ( .ip1(n9816), .ip2(\cache_data_B[7][36] ), .s(n9805), .op(
        n5428) );
  mux2_1 U12506 ( .ip1(n9817), .ip2(\cache_data_B[7][37] ), .s(n9805), .op(
        n5427) );
  mux2_1 U12507 ( .ip1(n9818), .ip2(\cache_data_B[7][38] ), .s(n9805), .op(
        n5426) );
  mux2_1 U12508 ( .ip1(n9819), .ip2(\cache_data_B[7][39] ), .s(n9805), .op(
        n5425) );
  mux2_1 U12509 ( .ip1(n9820), .ip2(\cache_data_B[7][40] ), .s(n9805), .op(
        n5424) );
  mux2_1 U12510 ( .ip1(n9821), .ip2(\cache_data_B[7][41] ), .s(n9805), .op(
        n5423) );
  buf_1 U12511 ( .ip(n9805), .op(n9806) );
  mux2_1 U12512 ( .ip1(n9822), .ip2(\cache_data_B[7][42] ), .s(n9806), .op(
        n5422) );
  mux2_1 U12513 ( .ip1(n9823), .ip2(\cache_data_B[7][43] ), .s(n9805), .op(
        n5421) );
  mux2_1 U12514 ( .ip1(n9824), .ip2(\cache_data_B[7][44] ), .s(n9805), .op(
        n5420) );
  mux2_1 U12515 ( .ip1(n9825), .ip2(\cache_data_B[7][45] ), .s(n9805), .op(
        n5419) );
  mux2_1 U12516 ( .ip1(n9826), .ip2(\cache_data_B[7][46] ), .s(n9805), .op(
        n5418) );
  mux2_1 U12517 ( .ip1(n9827), .ip2(\cache_data_B[7][47] ), .s(n9805), .op(
        n5417) );
  mux2_1 U12518 ( .ip1(n9828), .ip2(\cache_data_B[7][48] ), .s(n9806), .op(
        n5416) );
  mux2_1 U12519 ( .ip1(n9829), .ip2(\cache_data_B[7][49] ), .s(n9806), .op(
        n5415) );
  mux2_1 U12520 ( .ip1(n9830), .ip2(\cache_data_B[7][50] ), .s(n9806), .op(
        n5414) );
  mux2_1 U12521 ( .ip1(n9831), .ip2(\cache_data_B[7][51] ), .s(n9805), .op(
        n5413) );
  mux2_1 U12522 ( .ip1(n9832), .ip2(\cache_data_B[7][52] ), .s(n9805), .op(
        n5412) );
  mux2_1 U12523 ( .ip1(n9833), .ip2(\cache_data_B[7][53] ), .s(n9805), .op(
        n5411) );
  mux2_1 U12524 ( .ip1(n9835), .ip2(\cache_data_B[7][54] ), .s(n9805), .op(
        n5410) );
  mux2_1 U12525 ( .ip1(n9836), .ip2(\cache_data_B[7][55] ), .s(n9805), .op(
        n5409) );
  mux2_1 U12526 ( .ip1(n9837), .ip2(\cache_data_B[7][56] ), .s(n9805), .op(
        n5408) );
  mux2_1 U12527 ( .ip1(n9838), .ip2(\cache_data_B[7][57] ), .s(n9806), .op(
        n5407) );
  mux2_1 U12528 ( .ip1(n9839), .ip2(\cache_data_B[7][58] ), .s(n9806), .op(
        n5406) );
  mux2_1 U12529 ( .ip1(n9840), .ip2(\cache_data_B[7][59] ), .s(n9806), .op(
        n5405) );
  mux2_1 U12530 ( .ip1(n9841), .ip2(\cache_data_B[7][60] ), .s(n9806), .op(
        n5404) );
  mux2_1 U12531 ( .ip1(n9842), .ip2(\cache_data_B[7][61] ), .s(n9806), .op(
        n5403) );
  mux2_1 U12532 ( .ip1(n9843), .ip2(\cache_data_B[7][62] ), .s(n9806), .op(
        n5402) );
  mux2_1 U12533 ( .ip1(n9845), .ip2(\cache_data_B[7][63] ), .s(n9806), .op(
        n5401) );
  nand2_1 U12534 ( .ip1(n9811), .ip2(n9807), .op(n9808) );
  mux2_1 U12535 ( .ip1(n9831), .ip2(\cache_data_B[7][83] ), .s(n9808), .op(
        n5400) );
  mux2_1 U12536 ( .ip1(n9832), .ip2(\cache_data_B[7][84] ), .s(n9808), .op(
        n5399) );
  mux2_1 U12537 ( .ip1(n9833), .ip2(\cache_data_B[7][85] ), .s(n9808), .op(
        n5398) );
  mux2_1 U12538 ( .ip1(n9835), .ip2(\cache_data_B[7][86] ), .s(n9808), .op(
        n5397) );
  mux2_1 U12539 ( .ip1(n9836), .ip2(\cache_data_B[7][87] ), .s(n9808), .op(
        n5396) );
  mux2_1 U12540 ( .ip1(n9837), .ip2(\cache_data_B[7][88] ), .s(n9808), .op(
        n5395) );
  mux2_1 U12541 ( .ip1(n9838), .ip2(\cache_data_B[7][89] ), .s(n9808), .op(
        n5394) );
  mux2_1 U12542 ( .ip1(n9839), .ip2(\cache_data_B[7][90] ), .s(n9808), .op(
        n5393) );
  mux2_1 U12543 ( .ip1(n9840), .ip2(\cache_data_B[7][91] ), .s(n9808), .op(
        n5392) );
  mux2_1 U12544 ( .ip1(n9841), .ip2(\cache_data_B[7][92] ), .s(n9808), .op(
        n5391) );
  mux2_1 U12545 ( .ip1(n9842), .ip2(\cache_data_B[7][93] ), .s(n9808), .op(
        n5390) );
  mux2_1 U12546 ( .ip1(n9843), .ip2(\cache_data_B[7][94] ), .s(n9808), .op(
        n5389) );
  mux2_1 U12547 ( .ip1(n9845), .ip2(\cache_data_B[7][95] ), .s(n9808), .op(
        n5388) );
  mux2_1 U12548 ( .ip1(n9812), .ip2(\cache_data_B[7][64] ), .s(n9808), .op(
        n5387) );
  mux2_1 U12549 ( .ip1(n9813), .ip2(\cache_data_B[7][65] ), .s(n9808), .op(
        n5386) );
  mux2_1 U12550 ( .ip1(n9814), .ip2(\cache_data_B[7][66] ), .s(n9808), .op(
        n5385) );
  mux2_1 U12551 ( .ip1(n9815), .ip2(\cache_data_B[7][67] ), .s(n9808), .op(
        n5384) );
  mux2_1 U12552 ( .ip1(n9816), .ip2(\cache_data_B[7][68] ), .s(n9808), .op(
        n5383) );
  mux2_1 U12553 ( .ip1(n9817), .ip2(\cache_data_B[7][69] ), .s(n9808), .op(
        n5382) );
  buf_1 U12554 ( .ip(n9808), .op(n9809) );
  mux2_1 U12555 ( .ip1(n9818), .ip2(\cache_data_B[7][70] ), .s(n9809), .op(
        n5381) );
  mux2_1 U12556 ( .ip1(n9819), .ip2(\cache_data_B[7][71] ), .s(n9809), .op(
        n5380) );
  mux2_1 U12557 ( .ip1(n9820), .ip2(\cache_data_B[7][72] ), .s(n9809), .op(
        n5379) );
  mux2_1 U12558 ( .ip1(n9821), .ip2(\cache_data_B[7][73] ), .s(n9809), .op(
        n5378) );
  mux2_1 U12559 ( .ip1(n9822), .ip2(\cache_data_B[7][74] ), .s(n9809), .op(
        n5377) );
  mux2_1 U12560 ( .ip1(n9823), .ip2(\cache_data_B[7][75] ), .s(n9808), .op(
        n5376) );
  mux2_1 U12561 ( .ip1(n9824), .ip2(\cache_data_B[7][76] ), .s(n9808), .op(
        n5375) );
  mux2_1 U12562 ( .ip1(n9825), .ip2(\cache_data_B[7][77] ), .s(n9809), .op(
        n5374) );
  mux2_1 U12563 ( .ip1(n9826), .ip2(\cache_data_B[7][78] ), .s(n9809), .op(
        n5373) );
  mux2_1 U12564 ( .ip1(n9827), .ip2(\cache_data_B[7][79] ), .s(n9809), .op(
        n5372) );
  mux2_1 U12565 ( .ip1(n9828), .ip2(\cache_data_B[7][80] ), .s(n9809), .op(
        n5371) );
  mux2_1 U12566 ( .ip1(n9829), .ip2(\cache_data_B[7][81] ), .s(n9809), .op(
        n5370) );
  mux2_1 U12567 ( .ip1(n9830), .ip2(\cache_data_B[7][82] ), .s(n9809), .op(
        n5369) );
  nand2_1 U12568 ( .ip1(n9811), .ip2(n9810), .op(n9834) );
  mux2_1 U12569 ( .ip1(n9812), .ip2(\cache_data_B[7][96] ), .s(n9834), .op(
        n5368) );
  mux2_1 U12570 ( .ip1(n9813), .ip2(\cache_data_B[7][97] ), .s(n9834), .op(
        n5367) );
  mux2_1 U12571 ( .ip1(n9814), .ip2(\cache_data_B[7][98] ), .s(n9834), .op(
        n5366) );
  mux2_1 U12572 ( .ip1(n9815), .ip2(\cache_data_B[7][99] ), .s(n9834), .op(
        n5365) );
  mux2_1 U12573 ( .ip1(n9816), .ip2(\cache_data_B[7][100] ), .s(n9834), .op(
        n5364) );
  mux2_1 U12574 ( .ip1(n9817), .ip2(\cache_data_B[7][101] ), .s(n9834), .op(
        n5363) );
  mux2_1 U12575 ( .ip1(n9818), .ip2(\cache_data_B[7][102] ), .s(n9834), .op(
        n5362) );
  mux2_1 U12576 ( .ip1(n9819), .ip2(\cache_data_B[7][103] ), .s(n9834), .op(
        n5361) );
  mux2_1 U12577 ( .ip1(n9820), .ip2(\cache_data_B[7][104] ), .s(n9834), .op(
        n5360) );
  mux2_1 U12578 ( .ip1(n9821), .ip2(\cache_data_B[7][105] ), .s(n9834), .op(
        n5359) );
  mux2_1 U12579 ( .ip1(n9822), .ip2(\cache_data_B[7][106] ), .s(n9834), .op(
        n5358) );
  buf_1 U12580 ( .ip(n9834), .op(n9844) );
  mux2_1 U12581 ( .ip1(n9823), .ip2(\cache_data_B[7][107] ), .s(n9844), .op(
        n5357) );
  mux2_1 U12582 ( .ip1(n9824), .ip2(\cache_data_B[7][108] ), .s(n9834), .op(
        n5356) );
  mux2_1 U12583 ( .ip1(n9825), .ip2(\cache_data_B[7][109] ), .s(n9834), .op(
        n5355) );
  mux2_1 U12584 ( .ip1(n9826), .ip2(\cache_data_B[7][110] ), .s(n9834), .op(
        n5354) );
  mux2_1 U12585 ( .ip1(n9827), .ip2(\cache_data_B[7][111] ), .s(n9834), .op(
        n5353) );
  mux2_1 U12586 ( .ip1(n9828), .ip2(\cache_data_B[7][112] ), .s(n9834), .op(
        n5352) );
  mux2_1 U12587 ( .ip1(n9829), .ip2(\cache_data_B[7][113] ), .s(n9834), .op(
        n5351) );
  mux2_1 U12588 ( .ip1(n9830), .ip2(\cache_data_B[7][114] ), .s(n9834), .op(
        n5350) );
  mux2_1 U12589 ( .ip1(n9831), .ip2(\cache_data_B[7][115] ), .s(n9834), .op(
        n5349) );
  mux2_1 U12590 ( .ip1(n9832), .ip2(\cache_data_B[7][116] ), .s(n9844), .op(
        n5348) );
  mux2_1 U12591 ( .ip1(n9833), .ip2(\cache_data_B[7][117] ), .s(n9834), .op(
        n5347) );
  mux2_1 U12592 ( .ip1(n9835), .ip2(\cache_data_B[7][118] ), .s(n9834), .op(
        n5346) );
  mux2_1 U12593 ( .ip1(n9836), .ip2(\cache_data_B[7][119] ), .s(n9844), .op(
        n5345) );
  mux2_1 U12594 ( .ip1(n9837), .ip2(\cache_data_B[7][120] ), .s(n9844), .op(
        n5344) );
  mux2_1 U12595 ( .ip1(n9838), .ip2(\cache_data_B[7][121] ), .s(n9844), .op(
        n5343) );
  mux2_1 U12596 ( .ip1(n9839), .ip2(\cache_data_B[7][122] ), .s(n9844), .op(
        n5342) );
  mux2_1 U12597 ( .ip1(n9840), .ip2(\cache_data_B[7][123] ), .s(n9844), .op(
        n5341) );
  mux2_1 U12598 ( .ip1(n9841), .ip2(\cache_data_B[7][124] ), .s(n9844), .op(
        n5340) );
  mux2_1 U12599 ( .ip1(n9842), .ip2(\cache_data_B[7][125] ), .s(n9844), .op(
        n5339) );
  mux2_1 U12600 ( .ip1(n9843), .ip2(\cache_data_B[7][126] ), .s(n9844), .op(
        n5338) );
  mux2_1 U12601 ( .ip1(n9845), .ip2(\cache_data_B[7][127] ), .s(n9844), .op(
        n5337) );
  nand2_1 U12602 ( .ip1(n9846), .ip2(n9885), .op(n9848) );
  nand2_1 U12603 ( .ip1(n9848), .ip2(n9847), .op(n9856) );
  nand2_1 U12604 ( .ip1(n12370), .ip2(n9856), .op(n9849) );
  mux2_1 U12605 ( .ip1(n13294), .ip2(cache_dirty_B[0]), .s(n9849), .op(n5336)
         );
  nand2_1 U12606 ( .ip1(n10166), .ip2(n9856), .op(n9850) );
  mux2_1 U12607 ( .ip1(n13294), .ip2(cache_dirty_B[1]), .s(n9850), .op(n5335)
         );
  nand2_1 U12608 ( .ip1(n10426), .ip2(n9856), .op(n9851) );
  mux2_1 U12609 ( .ip1(n13294), .ip2(cache_dirty_B[2]), .s(n9851), .op(n5334)
         );
  nand2_1 U12610 ( .ip1(n11535), .ip2(n9856), .op(n9852) );
  mux2_1 U12611 ( .ip1(n13294), .ip2(cache_dirty_B[3]), .s(n9852), .op(n5333)
         );
  nand2_1 U12612 ( .ip1(n12054), .ip2(n9856), .op(n9853) );
  mux2_1 U12613 ( .ip1(n13294), .ip2(cache_dirty_B[4]), .s(n9853), .op(n5332)
         );
  nand2_1 U12614 ( .ip1(n11280), .ip2(n9856), .op(n9854) );
  mux2_1 U12615 ( .ip1(n13294), .ip2(cache_dirty_B[5]), .s(n9854), .op(n5331)
         );
  nand2_1 U12616 ( .ip1(n12458), .ip2(n9856), .op(n9855) );
  mux2_1 U12617 ( .ip1(n13294), .ip2(cache_dirty_B[6]), .s(n9855), .op(n5330)
         );
  nand2_1 U12618 ( .ip1(n10575), .ip2(n9856), .op(n9857) );
  mux2_1 U12619 ( .ip1(n9872), .ip2(cache_dirty_B[7]), .s(n9857), .op(n5329)
         );
  nor2_1 U12620 ( .ip1(n9859), .ip2(n9858), .op(n9874) );
  nor2_1 U12621 ( .ip1(n9874), .ip2(n9860), .op(n9861) );
  mux2_1 U12622 ( .ip1(cache_dirty_A[0]), .ip2(n9872), .s(n9861), .op(n5328)
         );
  nor2_1 U12623 ( .ip1(n9874), .ip2(n9862), .op(n9863) );
  mux2_1 U12624 ( .ip1(cache_dirty_A[1]), .ip2(n9872), .s(n9863), .op(n5327)
         );
  nor2_1 U12625 ( .ip1(n9874), .ip2(n9864), .op(n9865) );
  mux2_1 U12626 ( .ip1(cache_dirty_A[2]), .ip2(n13294), .s(n9865), .op(n5326)
         );
  nor2_1 U12627 ( .ip1(n9874), .ip2(n9866), .op(n9867) );
  mux2_1 U12628 ( .ip1(cache_dirty_A[3]), .ip2(n13294), .s(n9867), .op(n5325)
         );
  nor2_1 U12629 ( .ip1(n9874), .ip2(n9868), .op(n9869) );
  mux2_1 U12630 ( .ip1(cache_dirty_A[4]), .ip2(n13294), .s(n9869), .op(n5324)
         );
  nor2_1 U12631 ( .ip1(n9874), .ip2(n9870), .op(n9871) );
  mux2_1 U12632 ( .ip1(cache_dirty_A[5]), .ip2(n9872), .s(n9871), .op(n5323)
         );
  nor2_1 U12633 ( .ip1(n9874), .ip2(n9762), .op(n9873) );
  mux2_1 U12634 ( .ip1(cache_dirty_A[6]), .ip2(n13294), .s(n9873), .op(n5322)
         );
  nor2_1 U12635 ( .ip1(n9874), .ip2(n9769), .op(n9875) );
  mux2_1 U12636 ( .ip1(cache_dirty_A[7]), .ip2(n13294), .s(n9875), .op(n5321)
         );
  nor2_1 U12637 ( .ip1(n9885), .ip2(n9924), .op(n12550) );
  nand2_1 U12638 ( .ip1(\cache_data_A[7][0] ), .ip2(n12552), .op(n9884) );
  and2_1 U12639 ( .ip1(n11946), .ip2(\cache_data_A[1][0] ), .op(n9881) );
  nand2_1 U12640 ( .ip1(n12458), .ip2(\cache_data_A[6][0] ), .op(n9879) );
  nand2_1 U12641 ( .ip1(n11535), .ip2(\cache_data_A[3][0] ), .op(n9878) );
  nand2_1 U12642 ( .ip1(n11280), .ip2(\cache_data_A[5][0] ), .op(n9877) );
  nand2_1 U12643 ( .ip1(n12370), .ip2(\cache_data_A[0][0] ), .op(n9876) );
  nand4_1 U12644 ( .ip1(n9879), .ip2(n9878), .ip3(n9877), .ip4(n9876), .op(
        n9880) );
  not_ab_or_c_or_d U12645 ( .ip1(\cache_data_A[2][0] ), .ip2(n12475), .ip3(
        n9881), .ip4(n9880), .op(n9883) );
  nand2_1 U12646 ( .ip1(n12476), .ip2(\cache_data_A[4][0] ), .op(n9882) );
  nand3_1 U12647 ( .ip1(n9884), .ip2(n9883), .ip3(n9882), .op(n12605) );
  nand2_1 U12648 ( .ip1(n12550), .ip2(n12605), .op(n9961) );
  and2_1 U12649 ( .ip1(n9885), .ip2(n9905), .op(n12580) );
  nand2_1 U12650 ( .ip1(\cache_data_B[4][64] ), .ip2(n12194), .op(n9894) );
  and2_1 U12651 ( .ip1(n12429), .ip2(\cache_data_B[6][64] ), .op(n9891) );
  nand2_1 U12652 ( .ip1(n12370), .ip2(\cache_data_B[0][64] ), .op(n9889) );
  nand2_1 U12653 ( .ip1(n11535), .ip2(\cache_data_B[3][64] ), .op(n9888) );
  nand2_1 U12654 ( .ip1(n10426), .ip2(\cache_data_B[2][64] ), .op(n9887) );
  nand2_1 U12655 ( .ip1(n11280), .ip2(\cache_data_B[5][64] ), .op(n9886) );
  nand4_1 U12656 ( .ip1(n9889), .ip2(n9888), .ip3(n9887), .ip4(n9886), .op(
        n9890) );
  not_ab_or_c_or_d U12657 ( .ip1(\cache_data_B[7][64] ), .ip2(n12278), .ip3(
        n9891), .ip4(n9890), .op(n9893) );
  nand2_1 U12658 ( .ip1(n10166), .ip2(\cache_data_B[1][64] ), .op(n9892) );
  nand3_1 U12659 ( .ip1(n9894), .ip2(n9893), .ip3(n9892), .op(n12603) );
  nand2_1 U12660 ( .ip1(n10575), .ip2(\cache_data_A[7][64] ), .op(n9898) );
  nand2_1 U12661 ( .ip1(n10426), .ip2(\cache_data_A[2][64] ), .op(n9897) );
  nand2_1 U12662 ( .ip1(n11535), .ip2(\cache_data_A[3][64] ), .op(n9896) );
  nand2_1 U12663 ( .ip1(n11324), .ip2(\cache_data_A[4][64] ), .op(n9895) );
  nand4_1 U12664 ( .ip1(n9898), .ip2(n9897), .ip3(n9896), .ip4(n9895), .op(
        n9904) );
  nand2_1 U12665 ( .ip1(n11280), .ip2(\cache_data_A[5][64] ), .op(n9902) );
  nand2_1 U12666 ( .ip1(\cache_data_A[0][64] ), .ip2(n12204), .op(n9901) );
  nand2_1 U12667 ( .ip1(n10166), .ip2(\cache_data_A[1][64] ), .op(n9900) );
  nand2_1 U12668 ( .ip1(n12458), .ip2(\cache_data_A[6][64] ), .op(n9899) );
  nand4_1 U12669 ( .ip1(n9902), .ip2(n9901), .ip3(n9900), .ip4(n9899), .op(
        n9903) );
  nor2_1 U12670 ( .ip1(n9904), .ip2(n9903), .op(n12602) );
  nand2_1 U12671 ( .ip1(n9905), .ip2(n9925), .op(n12529) );
  nor2_1 U12672 ( .ip1(n12602), .ip2(n12529), .op(n9949) );
  nand2_1 U12673 ( .ip1(\cache_data_A[7][32] ), .ip2(n12552), .op(n9914) );
  and2_1 U12674 ( .ip1(n12147), .ip2(\cache_data_A[1][32] ), .op(n9911) );
  nand2_1 U12675 ( .ip1(n11280), .ip2(\cache_data_A[5][32] ), .op(n9909) );
  nand2_1 U12676 ( .ip1(n12584), .ip2(\cache_data_A[4][32] ), .op(n9908) );
  nand2_1 U12677 ( .ip1(n12458), .ip2(\cache_data_A[6][32] ), .op(n9907) );
  nand2_1 U12678 ( .ip1(n10426), .ip2(\cache_data_A[2][32] ), .op(n9906) );
  nand4_1 U12679 ( .ip1(n9909), .ip2(n9908), .ip3(n9907), .ip4(n9906), .op(
        n9910) );
  not_ab_or_c_or_d U12680 ( .ip1(\cache_data_A[0][32] ), .ip2(n12297), .ip3(
        n9911), .ip4(n9910), .op(n9913) );
  nand2_1 U12681 ( .ip1(n11535), .ip2(\cache_data_A[3][32] ), .op(n9912) );
  nand3_1 U12682 ( .ip1(n9914), .ip2(n9913), .ip3(n9912), .op(n12604) );
  nand2_1 U12683 ( .ip1(n12595), .ip2(n12604), .op(n9947) );
  nand2_1 U12684 ( .ip1(n10702), .ip2(\cache_data_B[7][32] ), .op(n9923) );
  and2_1 U12685 ( .ip1(n11780), .ip2(\cache_data_B[6][32] ), .op(n9920) );
  nand2_1 U12686 ( .ip1(n11156), .ip2(\cache_data_B[4][32] ), .op(n9918) );
  nand2_1 U12687 ( .ip1(n10426), .ip2(\cache_data_B[2][32] ), .op(n9917) );
  nand2_1 U12688 ( .ip1(n11535), .ip2(\cache_data_B[3][32] ), .op(n9916) );
  nand2_1 U12689 ( .ip1(n10166), .ip2(\cache_data_B[1][32] ), .op(n9915) );
  nand4_1 U12690 ( .ip1(n9918), .ip2(n9917), .ip3(n9916), .ip4(n9915), .op(
        n9919) );
  not_ab_or_c_or_d U12691 ( .ip1(\cache_data_B[0][32] ), .ip2(n12357), .ip3(
        n9920), .ip4(n9919), .op(n9922) );
  nand2_1 U12692 ( .ip1(n11280), .ip2(\cache_data_B[5][32] ), .op(n9921) );
  nand3_1 U12693 ( .ip1(n9923), .ip2(n9922), .ip3(n9921), .op(n12614) );
  nand2_1 U12694 ( .ip1(n12563), .ip2(n12614), .op(n9946) );
  nor2_1 U12695 ( .ip1(n9925), .ip2(n9924), .op(n12539) );
  nand2_1 U12696 ( .ip1(\cache_data_B[6][0] ), .ip2(n12371), .op(n9934) );
  and2_1 U12697 ( .ip1(n12486), .ip2(\cache_data_B[2][0] ), .op(n9931) );
  nand2_1 U12698 ( .ip1(n12278), .ip2(\cache_data_B[7][0] ), .op(n9929) );
  nand2_1 U12699 ( .ip1(n12054), .ip2(\cache_data_B[4][0] ), .op(n9928) );
  nand2_1 U12700 ( .ip1(n11280), .ip2(\cache_data_B[5][0] ), .op(n9927) );
  nand2_1 U12701 ( .ip1(n10166), .ip2(\cache_data_B[1][0] ), .op(n9926) );
  nand4_1 U12702 ( .ip1(n9929), .ip2(n9928), .ip3(n9927), .ip4(n9926), .op(
        n9930) );
  not_ab_or_c_or_d U12703 ( .ip1(\cache_data_B[0][0] ), .ip2(n12357), .ip3(
        n9931), .ip4(n9930), .op(n9933) );
  nand2_1 U12704 ( .ip1(n11535), .ip2(\cache_data_B[3][0] ), .op(n9932) );
  nand3_1 U12705 ( .ip1(n9934), .ip2(n9933), .ip3(n9932), .op(n12613) );
  nand2_1 U12706 ( .ip1(n12539), .ip2(n12613), .op(n9945) );
  nand2_1 U12707 ( .ip1(n11535), .ip2(\cache_data_A[3][96] ), .op(n9943) );
  and2_1 U12708 ( .ip1(n12147), .ip2(\cache_data_A[1][96] ), .op(n9940) );
  nand2_1 U12709 ( .ip1(n11156), .ip2(\cache_data_A[4][96] ), .op(n9938) );
  nand2_1 U12710 ( .ip1(n12468), .ip2(\cache_data_A[7][96] ), .op(n9937) );
  nand2_1 U12711 ( .ip1(n12370), .ip2(\cache_data_A[0][96] ), .op(n9936) );
  nand2_1 U12712 ( .ip1(n12458), .ip2(\cache_data_A[6][96] ), .op(n9935) );
  nand4_1 U12713 ( .ip1(n9938), .ip2(n9937), .ip3(n9936), .ip4(n9935), .op(
        n9939) );
  not_ab_or_c_or_d U12714 ( .ip1(\cache_data_A[2][96] ), .ip2(n12475), .ip3(
        n9940), .ip4(n9939), .op(n9942) );
  nand2_1 U12715 ( .ip1(n11280), .ip2(\cache_data_A[5][96] ), .op(n9941) );
  nand3_1 U12716 ( .ip1(n9943), .ip2(n9942), .ip3(n9941), .op(n12601) );
  nand2_1 U12717 ( .ip1(n12509), .ip2(n12601), .op(n9944) );
  nand4_1 U12718 ( .ip1(n9947), .ip2(n9946), .ip3(n9945), .ip4(n9944), .op(
        n9948) );
  not_ab_or_c_or_d U12719 ( .ip1(n12580), .ip2(n12603), .ip3(n9949), .ip4(
        n9948), .op(n9960) );
  nand2_1 U12720 ( .ip1(\cache_data_B[0][96] ), .ip2(n12204), .op(n9958) );
  and2_1 U12721 ( .ip1(n12582), .ip2(\cache_data_B[5][96] ), .op(n9955) );
  nand2_1 U12722 ( .ip1(n12458), .ip2(\cache_data_B[6][96] ), .op(n9953) );
  nand2_1 U12723 ( .ip1(n10166), .ip2(\cache_data_B[1][96] ), .op(n9952) );
  nand2_1 U12724 ( .ip1(n10575), .ip2(\cache_data_B[7][96] ), .op(n9951) );
  nand2_1 U12725 ( .ip1(n10426), .ip2(\cache_data_B[2][96] ), .op(n9950) );
  nand4_1 U12726 ( .ip1(n9953), .ip2(n9952), .ip3(n9951), .ip4(n9950), .op(
        n9954) );
  not_ab_or_c_or_d U12727 ( .ip1(\cache_data_B[4][96] ), .ip2(n12476), .ip3(
        n9955), .ip4(n9954), .op(n9957) );
  nand2_1 U12728 ( .ip1(n12096), .ip2(\cache_data_B[3][96] ), .op(n9956) );
  nand3_1 U12729 ( .ip1(n9958), .ip2(n9957), .ip3(n9956), .op(n12606) );
  nand2_1 U12730 ( .ip1(n12573), .ip2(n12606), .op(n9959) );
  nand3_1 U12731 ( .ip1(n9961), .ip2(n9960), .ip3(n9959), .op(n9962) );
  mux2_1 U12732 ( .ip1(N4204), .ip2(n9962), .s(n10378), .op(n5320) );
  nand2_1 U12733 ( .ip1(n10426), .ip2(\cache_data_A[2][33] ), .op(n9971) );
  and2_1 U12734 ( .ip1(n10686), .ip2(\cache_data_A[1][33] ), .op(n9968) );
  nand2_1 U12735 ( .ip1(n12584), .ip2(\cache_data_A[4][33] ), .op(n9966) );
  nand2_1 U12736 ( .ip1(n12458), .ip2(\cache_data_A[6][33] ), .op(n9965) );
  nand2_1 U12737 ( .ip1(n12370), .ip2(\cache_data_A[0][33] ), .op(n9964) );
  nand2_1 U12738 ( .ip1(n11280), .ip2(\cache_data_A[5][33] ), .op(n9963) );
  nand4_1 U12739 ( .ip1(n9966), .ip2(n9965), .ip3(n9964), .ip4(n9963), .op(
        n9967) );
  not_ab_or_c_or_d U12740 ( .ip1(\cache_data_A[3][33] ), .ip2(n11535), .ip3(
        n9968), .ip4(n9967), .op(n9970) );
  nand2_1 U12741 ( .ip1(n11057), .ip2(\cache_data_A[7][33] ), .op(n9969) );
  nand3_1 U12742 ( .ip1(n9971), .ip2(n9970), .ip3(n9969), .op(n12622) );
  nand2_1 U12743 ( .ip1(n12595), .ip2(n12622), .op(n10044) );
  nand2_1 U12744 ( .ip1(\cache_data_B[1][97] ), .ip2(n11724), .op(n9980) );
  and2_1 U12745 ( .ip1(n12486), .ip2(\cache_data_B[2][97] ), .op(n9977) );
  nand2_1 U12746 ( .ip1(n12458), .ip2(\cache_data_B[6][97] ), .op(n9975) );
  nand2_1 U12747 ( .ip1(n12559), .ip2(\cache_data_B[3][97] ), .op(n9974) );
  nand2_1 U12748 ( .ip1(n12054), .ip2(\cache_data_B[4][97] ), .op(n9973) );
  nand2_1 U12749 ( .ip1(n11057), .ip2(\cache_data_B[7][97] ), .op(n9972) );
  nand4_1 U12750 ( .ip1(n9975), .ip2(n9974), .ip3(n9973), .ip4(n9972), .op(
        n9976) );
  not_ab_or_c_or_d U12751 ( .ip1(\cache_data_B[0][97] ), .ip2(n12357), .ip3(
        n9977), .ip4(n9976), .op(n9979) );
  nand2_1 U12752 ( .ip1(n11280), .ip2(\cache_data_B[5][97] ), .op(n9978) );
  nand3_1 U12753 ( .ip1(n9980), .ip2(n9979), .ip3(n9978), .op(n12624) );
  nand2_1 U12754 ( .ip1(n11280), .ip2(\cache_data_A[5][65] ), .op(n9984) );
  nand2_1 U12755 ( .ip1(n12096), .ip2(\cache_data_A[3][65] ), .op(n9983) );
  nand2_1 U12756 ( .ip1(n10702), .ip2(\cache_data_A[7][65] ), .op(n9982) );
  nand2_1 U12757 ( .ip1(n10426), .ip2(\cache_data_A[2][65] ), .op(n9981) );
  nand4_1 U12758 ( .ip1(n9984), .ip2(n9983), .ip3(n9982), .ip4(n9981), .op(
        n9990) );
  nand2_1 U12759 ( .ip1(n10166), .ip2(\cache_data_A[1][65] ), .op(n9988) );
  nand2_1 U12760 ( .ip1(n12370), .ip2(\cache_data_A[0][65] ), .op(n9987) );
  nand2_1 U12761 ( .ip1(n12054), .ip2(\cache_data_A[4][65] ), .op(n9986) );
  nand2_1 U12762 ( .ip1(n11780), .ip2(\cache_data_A[6][65] ), .op(n9985) );
  nand4_1 U12763 ( .ip1(n9988), .ip2(n9987), .ip3(n9986), .ip4(n9985), .op(
        n9989) );
  nor2_1 U12764 ( .ip1(n9990), .ip2(n9989), .op(n12621) );
  nor2_1 U12765 ( .ip1(n12621), .ip2(n12529), .op(n10032) );
  nand2_1 U12766 ( .ip1(n12096), .ip2(\cache_data_A[3][1] ), .op(n9999) );
  and2_1 U12767 ( .ip1(n12476), .ip2(\cache_data_A[4][1] ), .op(n9996) );
  nand2_1 U12768 ( .ip1(n12370), .ip2(\cache_data_A[0][1] ), .op(n9994) );
  nand2_1 U12769 ( .ip1(n11057), .ip2(\cache_data_A[7][1] ), .op(n9993) );
  nand2_1 U12770 ( .ip1(n10426), .ip2(\cache_data_A[2][1] ), .op(n9992) );
  nand2_1 U12771 ( .ip1(n11280), .ip2(\cache_data_A[5][1] ), .op(n9991) );
  nand4_1 U12772 ( .ip1(n9994), .ip2(n9993), .ip3(n9992), .ip4(n9991), .op(
        n9995) );
  not_ab_or_c_or_d U12773 ( .ip1(\cache_data_A[6][1] ), .ip2(n12337), .ip3(
        n9996), .ip4(n9995), .op(n9998) );
  nand2_1 U12774 ( .ip1(n10166), .ip2(\cache_data_A[1][1] ), .op(n9997) );
  nand3_1 U12775 ( .ip1(n9999), .ip2(n9998), .ip3(n9997), .op(n12623) );
  nand2_1 U12776 ( .ip1(n12550), .ip2(n12623), .op(n10030) );
  nand2_1 U12777 ( .ip1(\cache_data_B[6][33] ), .ip2(n12458), .op(n10008) );
  and2_1 U12778 ( .ip1(n12581), .ip2(\cache_data_B[7][33] ), .op(n10005) );
  nand2_1 U12779 ( .ip1(n11535), .ip2(\cache_data_B[3][33] ), .op(n10003) );
  nand2_1 U12780 ( .ip1(n12054), .ip2(\cache_data_B[4][33] ), .op(n10002) );
  nand2_1 U12781 ( .ip1(n10426), .ip2(\cache_data_B[2][33] ), .op(n10001) );
  nand2_1 U12782 ( .ip1(n10166), .ip2(\cache_data_B[1][33] ), .op(n10000) );
  nand4_1 U12783 ( .ip1(n10003), .ip2(n10002), .ip3(n10001), .ip4(n10000), 
        .op(n10004) );
  not_ab_or_c_or_d U12784 ( .ip1(\cache_data_B[0][33] ), .ip2(n12357), .ip3(
        n10005), .ip4(n10004), .op(n10007) );
  nand2_1 U12785 ( .ip1(n11280), .ip2(\cache_data_B[5][33] ), .op(n10006) );
  nand3_1 U12786 ( .ip1(n10008), .ip2(n10007), .ip3(n10006), .op(n12625) );
  nand2_1 U12787 ( .ip1(n12563), .ip2(n12625), .op(n10029) );
  nand2_1 U12788 ( .ip1(\cache_data_A[0][97] ), .ip2(n12204), .op(n10017) );
  and2_1 U12789 ( .ip1(n12147), .ip2(\cache_data_A[1][97] ), .op(n10014) );
  nand2_1 U12790 ( .ip1(n10426), .ip2(\cache_data_A[2][97] ), .op(n10012) );
  nand2_1 U12791 ( .ip1(n11780), .ip2(\cache_data_A[6][97] ), .op(n10011) );
  nand2_1 U12792 ( .ip1(n12054), .ip2(\cache_data_A[4][97] ), .op(n10010) );
  nand2_1 U12793 ( .ip1(n12581), .ip2(\cache_data_A[7][97] ), .op(n10009) );
  nand4_1 U12794 ( .ip1(n10012), .ip2(n10011), .ip3(n10010), .ip4(n10009), 
        .op(n10013) );
  not_ab_or_c_or_d U12795 ( .ip1(\cache_data_A[3][97] ), .ip2(n11535), .ip3(
        n10014), .ip4(n10013), .op(n10016) );
  nand2_1 U12796 ( .ip1(n11236), .ip2(\cache_data_A[5][97] ), .op(n10015) );
  nand3_1 U12797 ( .ip1(n10017), .ip2(n10016), .ip3(n10015), .op(n12620) );
  nand2_1 U12798 ( .ip1(n12509), .ip2(n12620), .op(n10028) );
  nand2_1 U12799 ( .ip1(n10426), .ip2(\cache_data_B[2][65] ), .op(n10026) );
  and2_1 U12800 ( .ip1(n12476), .ip2(\cache_data_B[4][65] ), .op(n10023) );
  nand2_1 U12801 ( .ip1(n12370), .ip2(\cache_data_B[0][65] ), .op(n10021) );
  nand2_1 U12802 ( .ip1(n10166), .ip2(\cache_data_B[1][65] ), .op(n10020) );
  nand2_1 U12803 ( .ip1(n11780), .ip2(\cache_data_B[6][65] ), .op(n10019) );
  nand2_1 U12804 ( .ip1(n10702), .ip2(\cache_data_B[7][65] ), .op(n10018) );
  nand4_1 U12805 ( .ip1(n10021), .ip2(n10020), .ip3(n10019), .ip4(n10018), 
        .op(n10022) );
  not_ab_or_c_or_d U12806 ( .ip1(\cache_data_B[3][65] ), .ip2(n11535), .ip3(
        n10023), .ip4(n10022), .op(n10025) );
  nand2_1 U12807 ( .ip1(n11236), .ip2(\cache_data_B[5][65] ), .op(n10024) );
  nand3_1 U12808 ( .ip1(n10026), .ip2(n10025), .ip3(n10024), .op(n12632) );
  nand2_1 U12809 ( .ip1(n12580), .ip2(n12632), .op(n10027) );
  nand4_1 U12810 ( .ip1(n10030), .ip2(n10029), .ip3(n10028), .ip4(n10027), 
        .op(n10031) );
  not_ab_or_c_or_d U12811 ( .ip1(n12573), .ip2(n12624), .ip3(n10032), .ip4(
        n10031), .op(n10043) );
  nand2_1 U12812 ( .ip1(n12370), .ip2(\cache_data_B[0][1] ), .op(n10041) );
  and2_1 U12813 ( .ip1(n12581), .ip2(\cache_data_B[7][1] ), .op(n10038) );
  nand2_1 U12814 ( .ip1(n11236), .ip2(\cache_data_B[5][1] ), .op(n10036) );
  nand2_1 U12815 ( .ip1(n11780), .ip2(\cache_data_B[6][1] ), .op(n10035) );
  nand2_1 U12816 ( .ip1(n11724), .ip2(\cache_data_B[1][1] ), .op(n10034) );
  nand2_1 U12817 ( .ip1(n12559), .ip2(\cache_data_B[3][1] ), .op(n10033) );
  nand4_1 U12818 ( .ip1(n10036), .ip2(n10035), .ip3(n10034), .ip4(n10033), 
        .op(n10037) );
  not_ab_or_c_or_d U12819 ( .ip1(n12546), .ip2(\cache_data_B[2][1] ), .ip3(
        n10038), .ip4(n10037), .op(n10040) );
  nand2_1 U12820 ( .ip1(n11324), .ip2(\cache_data_B[4][1] ), .op(n10039) );
  nand3_1 U12821 ( .ip1(n10041), .ip2(n10040), .ip3(n10039), .op(n12633) );
  nand2_1 U12822 ( .ip1(n12539), .ip2(n12633), .op(n10042) );
  nand3_1 U12823 ( .ip1(n10044), .ip2(n10043), .ip3(n10042), .op(n10045) );
  mux2_1 U12824 ( .ip1(N4201), .ip2(n10045), .s(n10378), .op(n5319) );
  nand2_1 U12825 ( .ip1(\cache_data_A[0][34] ), .ip2(n12204), .op(n10054) );
  and2_1 U12826 ( .ip1(n8060), .ip2(\cache_data_A[3][34] ), .op(n10051) );
  nand2_1 U12827 ( .ip1(n12371), .ip2(\cache_data_A[6][34] ), .op(n10049) );
  nand2_1 U12828 ( .ip1(n11724), .ip2(\cache_data_A[1][34] ), .op(n10048) );
  nand2_1 U12829 ( .ip1(n11236), .ip2(\cache_data_A[5][34] ), .op(n10047) );
  nand2_1 U12830 ( .ip1(n11324), .ip2(\cache_data_A[4][34] ), .op(n10046) );
  nand4_1 U12831 ( .ip1(n10049), .ip2(n10048), .ip3(n10047), .ip4(n10046), 
        .op(n10050) );
  not_ab_or_c_or_d U12832 ( .ip1(\cache_data_A[2][34] ), .ip2(n12546), .ip3(
        n10051), .ip4(n10050), .op(n10053) );
  nand2_1 U12833 ( .ip1(n12581), .ip2(\cache_data_A[7][34] ), .op(n10052) );
  nand3_1 U12834 ( .ip1(n10054), .ip2(n10053), .ip3(n10052), .op(n12651) );
  nand2_1 U12835 ( .ip1(n12595), .ip2(n12651), .op(n10127) );
  nand2_1 U12836 ( .ip1(n10426), .ip2(\cache_data_B[2][66] ), .op(n10063) );
  and2_1 U12837 ( .ip1(n12476), .ip2(\cache_data_B[4][66] ), .op(n10060) );
  nand2_1 U12838 ( .ip1(n10166), .ip2(\cache_data_B[1][66] ), .op(n10058) );
  nand2_1 U12839 ( .ip1(n12581), .ip2(\cache_data_B[7][66] ), .op(n10057) );
  nand2_1 U12840 ( .ip1(n11535), .ip2(\cache_data_B[3][66] ), .op(n10056) );
  nand2_1 U12841 ( .ip1(n12458), .ip2(\cache_data_B[6][66] ), .op(n10055) );
  nand4_1 U12842 ( .ip1(n10058), .ip2(n10057), .ip3(n10056), .ip4(n10055), 
        .op(n10059) );
  not_ab_or_c_or_d U12843 ( .ip1(n8452), .ip2(\cache_data_B[0][66] ), .ip3(
        n10060), .ip4(n10059), .op(n10062) );
  nand2_1 U12844 ( .ip1(n11236), .ip2(\cache_data_B[5][66] ), .op(n10061) );
  nand3_1 U12845 ( .ip1(n10063), .ip2(n10062), .ip3(n10061), .op(n12640) );
  nand2_1 U12846 ( .ip1(n12559), .ip2(\cache_data_A[3][66] ), .op(n10067) );
  nand2_1 U12847 ( .ip1(n12370), .ip2(\cache_data_A[0][66] ), .op(n10066) );
  nand2_1 U12848 ( .ip1(n10426), .ip2(\cache_data_A[2][66] ), .op(n10065) );
  nand2_1 U12849 ( .ip1(n12581), .ip2(\cache_data_A[7][66] ), .op(n10064) );
  nand4_1 U12850 ( .ip1(n10067), .ip2(n10066), .ip3(n10065), .ip4(n10064), 
        .op(n10073) );
  nand2_1 U12851 ( .ip1(n11780), .ip2(\cache_data_A[6][66] ), .op(n10071) );
  nand2_1 U12852 ( .ip1(n11724), .ip2(\cache_data_A[1][66] ), .op(n10070) );
  nand2_1 U12853 ( .ip1(n11324), .ip2(\cache_data_A[4][66] ), .op(n10069) );
  nand2_1 U12854 ( .ip1(n11236), .ip2(\cache_data_A[5][66] ), .op(n10068) );
  nand4_1 U12855 ( .ip1(n10071), .ip2(n10070), .ip3(n10069), .ip4(n10068), 
        .op(n10072) );
  nor2_1 U12856 ( .ip1(n10073), .ip2(n10072), .op(n12639) );
  nor2_1 U12857 ( .ip1(n12639), .ip2(n12529), .op(n10115) );
  nand2_1 U12858 ( .ip1(n12559), .ip2(\cache_data_A[3][98] ), .op(n10082) );
  and2_1 U12859 ( .ip1(n12320), .ip2(\cache_data_A[6][98] ), .op(n10079) );
  nand2_1 U12860 ( .ip1(n11324), .ip2(\cache_data_A[4][98] ), .op(n10077) );
  nand2_1 U12861 ( .ip1(n12581), .ip2(\cache_data_A[7][98] ), .op(n10076) );
  nand2_1 U12862 ( .ip1(n10166), .ip2(\cache_data_A[1][98] ), .op(n10075) );
  nand2_1 U12863 ( .ip1(n12370), .ip2(\cache_data_A[0][98] ), .op(n10074) );
  nand4_1 U12864 ( .ip1(n10077), .ip2(n10076), .ip3(n10075), .ip4(n10074), 
        .op(n10078) );
  not_ab_or_c_or_d U12865 ( .ip1(\cache_data_A[2][98] ), .ip2(n12546), .ip3(
        n10079), .ip4(n10078), .op(n10081) );
  nand2_1 U12866 ( .ip1(n11236), .ip2(\cache_data_A[5][98] ), .op(n10080) );
  nand3_1 U12867 ( .ip1(n10082), .ip2(n10081), .ip3(n10080), .op(n12650) );
  nand2_1 U12868 ( .ip1(n12509), .ip2(n12650), .op(n10113) );
  nand2_1 U12869 ( .ip1(n11071), .ip2(\cache_data_A[0][2] ), .op(n10091) );
  and2_1 U12870 ( .ip1(n12468), .ip2(\cache_data_A[7][2] ), .op(n10088) );
  nand2_1 U12871 ( .ip1(n11535), .ip2(\cache_data_A[3][2] ), .op(n10086) );
  nand2_1 U12872 ( .ip1(n12054), .ip2(\cache_data_A[4][2] ), .op(n10085) );
  nand2_1 U12873 ( .ip1(n12371), .ip2(\cache_data_A[6][2] ), .op(n10084) );
  nand2_1 U12874 ( .ip1(n11236), .ip2(\cache_data_A[5][2] ), .op(n10083) );
  nand4_1 U12875 ( .ip1(n10086), .ip2(n10085), .ip3(n10084), .ip4(n10083), 
        .op(n10087) );
  not_ab_or_c_or_d U12876 ( .ip1(\cache_data_A[2][2] ), .ip2(n12475), .ip3(
        n10088), .ip4(n10087), .op(n10090) );
  nand2_1 U12877 ( .ip1(n10166), .ip2(\cache_data_A[1][2] ), .op(n10089) );
  nand3_1 U12878 ( .ip1(n10091), .ip2(n10090), .ip3(n10089), .op(n12638) );
  nand2_1 U12879 ( .ip1(n12550), .ip2(n12638), .op(n10112) );
  nand2_1 U12880 ( .ip1(\cache_data_B[0][98] ), .ip2(n12204), .op(n10100) );
  and2_1 U12881 ( .ip1(n12396), .ip2(\cache_data_B[4][98] ), .op(n10097) );
  nand2_1 U12882 ( .ip1(n10426), .ip2(\cache_data_B[2][98] ), .op(n10095) );
  nand2_1 U12883 ( .ip1(n12581), .ip2(\cache_data_B[7][98] ), .op(n10094) );
  nand2_1 U12884 ( .ip1(n11236), .ip2(\cache_data_B[5][98] ), .op(n10093) );
  nand2_1 U12885 ( .ip1(n12096), .ip2(\cache_data_B[3][98] ), .op(n10092) );
  nand4_1 U12886 ( .ip1(n10095), .ip2(n10094), .ip3(n10093), .ip4(n10092), 
        .op(n10096) );
  not_ab_or_c_or_d U12887 ( .ip1(n12551), .ip2(\cache_data_B[6][98] ), .ip3(
        n10097), .ip4(n10096), .op(n10099) );
  nand2_1 U12888 ( .ip1(n11724), .ip2(\cache_data_B[1][98] ), .op(n10098) );
  nand3_1 U12889 ( .ip1(n10100), .ip2(n10099), .ip3(n10098), .op(n12642) );
  nand2_1 U12890 ( .ip1(n12573), .ip2(n12642), .op(n10111) );
  nand2_1 U12891 ( .ip1(\cache_data_B[0][34] ), .ip2(n12204), .op(n10109) );
  and2_1 U12892 ( .ip1(n12581), .ip2(\cache_data_B[7][34] ), .op(n10106) );
  nand2_1 U12893 ( .ip1(n12371), .ip2(\cache_data_B[6][34] ), .op(n10104) );
  nand2_1 U12894 ( .ip1(n10166), .ip2(\cache_data_B[1][34] ), .op(n10103) );
  nand2_1 U12895 ( .ip1(n12054), .ip2(\cache_data_B[4][34] ), .op(n10102) );
  nand2_1 U12896 ( .ip1(n11236), .ip2(\cache_data_B[5][34] ), .op(n10101) );
  nand4_1 U12897 ( .ip1(n10104), .ip2(n10103), .ip3(n10102), .ip4(n10101), 
        .op(n10105) );
  not_ab_or_c_or_d U12898 ( .ip1(\cache_data_B[2][34] ), .ip2(n12475), .ip3(
        n10106), .ip4(n10105), .op(n10108) );
  nand2_1 U12899 ( .ip1(n11535), .ip2(\cache_data_B[3][34] ), .op(n10107) );
  nand3_1 U12900 ( .ip1(n10109), .ip2(n10108), .ip3(n10107), .op(n12643) );
  nand2_1 U12901 ( .ip1(n12563), .ip2(n12643), .op(n10110) );
  nand4_1 U12902 ( .ip1(n10113), .ip2(n10112), .ip3(n10111), .ip4(n10110), 
        .op(n10114) );
  not_ab_or_c_or_d U12903 ( .ip1(n12580), .ip2(n12640), .ip3(n10115), .ip4(
        n10114), .op(n10126) );
  nand2_1 U12904 ( .ip1(n12468), .ip2(\cache_data_B[7][2] ), .op(n10124) );
  and2_1 U12905 ( .ip1(n12486), .ip2(\cache_data_B[2][2] ), .op(n10121) );
  nand2_1 U12906 ( .ip1(n11780), .ip2(\cache_data_B[6][2] ), .op(n10119) );
  nand2_1 U12907 ( .ip1(n11236), .ip2(\cache_data_B[5][2] ), .op(n10118) );
  nand2_1 U12908 ( .ip1(n11535), .ip2(\cache_data_B[3][2] ), .op(n10117) );
  nand2_1 U12909 ( .ip1(n10166), .ip2(\cache_data_B[1][2] ), .op(n10116) );
  nand4_1 U12910 ( .ip1(n10119), .ip2(n10118), .ip3(n10117), .ip4(n10116), 
        .op(n10120) );
  not_ab_or_c_or_d U12911 ( .ip1(\cache_data_B[0][2] ), .ip2(n12297), .ip3(
        n10121), .ip4(n10120), .op(n10123) );
  nand2_1 U12912 ( .ip1(n11324), .ip2(\cache_data_B[4][2] ), .op(n10122) );
  nand3_1 U12913 ( .ip1(n10124), .ip2(n10123), .ip3(n10122), .op(n12641) );
  nand2_1 U12914 ( .ip1(n12539), .ip2(n12641), .op(n10125) );
  nand3_1 U12915 ( .ip1(n10127), .ip2(n10126), .ip3(n10125), .op(n10128) );
  mux2_1 U12916 ( .ip1(N4198), .ip2(n10128), .s(n10378), .op(n5318) );
  nand2_1 U12917 ( .ip1(n12096), .ip2(\cache_data_B[3][67] ), .op(n10137) );
  and2_1 U12918 ( .ip1(n12396), .ip2(\cache_data_B[4][67] ), .op(n10134) );
  nand2_1 U12919 ( .ip1(n11296), .ip2(\cache_data_B[5][67] ), .op(n10132) );
  nand2_1 U12920 ( .ip1(n11780), .ip2(\cache_data_B[6][67] ), .op(n10131) );
  nand2_1 U12921 ( .ip1(n10426), .ip2(\cache_data_B[2][67] ), .op(n10130) );
  nand2_1 U12922 ( .ip1(n11071), .ip2(\cache_data_B[0][67] ), .op(n10129) );
  nand4_1 U12923 ( .ip1(n10132), .ip2(n10131), .ip3(n10130), .ip4(n10129), 
        .op(n10133) );
  not_ab_or_c_or_d U12924 ( .ip1(\cache_data_B[7][67] ), .ip2(n11057), .ip3(
        n10134), .ip4(n10133), .op(n10136) );
  nand2_1 U12925 ( .ip1(n11724), .ip2(\cache_data_B[1][67] ), .op(n10135) );
  nand3_1 U12926 ( .ip1(n10137), .ip2(n10136), .ip3(n10135), .op(n12661) );
  nand2_1 U12927 ( .ip1(n12580), .ip2(n12661), .op(n10211) );
  nand2_1 U12928 ( .ip1(\cache_data_B[6][3] ), .ip2(n12458), .op(n10146) );
  and2_1 U12929 ( .ip1(n12256), .ip2(\cache_data_B[5][3] ), .op(n10143) );
  nand2_1 U12930 ( .ip1(n10426), .ip2(\cache_data_B[2][3] ), .op(n10141) );
  nand2_1 U12931 ( .ip1(n11535), .ip2(\cache_data_B[3][3] ), .op(n10140) );
  nand2_1 U12932 ( .ip1(n10166), .ip2(\cache_data_B[1][3] ), .op(n10139) );
  nand2_1 U12933 ( .ip1(n11071), .ip2(\cache_data_B[0][3] ), .op(n10138) );
  nand4_1 U12934 ( .ip1(n10141), .ip2(n10140), .ip3(n10139), .ip4(n10138), 
        .op(n10142) );
  not_ab_or_c_or_d U12935 ( .ip1(\cache_data_B[7][3] ), .ip2(n12552), .ip3(
        n10143), .ip4(n10142), .op(n10145) );
  nand2_1 U12936 ( .ip1(n11156), .ip2(\cache_data_B[4][3] ), .op(n10144) );
  nand3_1 U12937 ( .ip1(n10146), .ip2(n10145), .ip3(n10144), .op(n12659) );
  nand2_1 U12938 ( .ip1(n10702), .ip2(\cache_data_A[7][67] ), .op(n10150) );
  nand2_1 U12939 ( .ip1(n11071), .ip2(\cache_data_A[0][67] ), .op(n10149) );
  nand2_1 U12940 ( .ip1(n12559), .ip2(\cache_data_A[3][67] ), .op(n10148) );
  nand2_1 U12941 ( .ip1(n10426), .ip2(\cache_data_A[2][67] ), .op(n10147) );
  nand4_1 U12942 ( .ip1(n10150), .ip2(n10149), .ip3(n10148), .ip4(n10147), 
        .op(n10156) );
  nand2_1 U12943 ( .ip1(n12320), .ip2(\cache_data_A[6][67] ), .op(n10154) );
  nand2_1 U12944 ( .ip1(n11236), .ip2(\cache_data_A[5][67] ), .op(n10153) );
  nand2_1 U12945 ( .ip1(n11724), .ip2(\cache_data_A[1][67] ), .op(n10152) );
  nand2_1 U12946 ( .ip1(n11156), .ip2(\cache_data_A[4][67] ), .op(n10151) );
  nand4_1 U12947 ( .ip1(n10154), .ip2(n10153), .ip3(n10152), .ip4(n10151), 
        .op(n10155) );
  nor2_1 U12948 ( .ip1(n10156), .ip2(n10155), .op(n12657) );
  nor2_1 U12949 ( .ip1(n12657), .ip2(n12529), .op(n10199) );
  nand2_1 U12950 ( .ip1(n12371), .ip2(\cache_data_A[6][3] ), .op(n10165) );
  and2_1 U12951 ( .ip1(n12396), .ip2(\cache_data_A[4][3] ), .op(n10162) );
  nand2_1 U12952 ( .ip1(n12468), .ip2(\cache_data_A[7][3] ), .op(n10160) );
  nand2_1 U12953 ( .ip1(n12559), .ip2(\cache_data_A[3][3] ), .op(n10159) );
  nand2_1 U12954 ( .ip1(n11296), .ip2(\cache_data_A[5][3] ), .op(n10158) );
  nand2_1 U12955 ( .ip1(n11071), .ip2(\cache_data_A[0][3] ), .op(n10157) );
  nand4_1 U12956 ( .ip1(n10160), .ip2(n10159), .ip3(n10158), .ip4(n10157), 
        .op(n10161) );
  not_ab_or_c_or_d U12957 ( .ip1(\cache_data_A[2][3] ), .ip2(n12546), .ip3(
        n10162), .ip4(n10161), .op(n10164) );
  nand2_1 U12958 ( .ip1(n11724), .ip2(\cache_data_A[1][3] ), .op(n10163) );
  nand3_1 U12959 ( .ip1(n10165), .ip2(n10164), .ip3(n10163), .op(n12668) );
  nand2_1 U12960 ( .ip1(n12550), .ip2(n12668), .op(n10197) );
  nand2_1 U12961 ( .ip1(\cache_data_B[3][35] ), .ip2(n12321), .op(n10175) );
  and2_1 U12962 ( .ip1(n11780), .ip2(\cache_data_B[6][35] ), .op(n10172) );
  nand2_1 U12963 ( .ip1(n11071), .ip2(\cache_data_B[0][35] ), .op(n10170) );
  nand2_1 U12964 ( .ip1(n10166), .ip2(\cache_data_B[1][35] ), .op(n10169) );
  nand2_1 U12965 ( .ip1(n10426), .ip2(\cache_data_B[2][35] ), .op(n10168) );
  nand2_1 U12966 ( .ip1(n12054), .ip2(\cache_data_B[4][35] ), .op(n10167) );
  nand4_1 U12967 ( .ip1(n10170), .ip2(n10169), .ip3(n10168), .ip4(n10167), 
        .op(n10171) );
  not_ab_or_c_or_d U12968 ( .ip1(n12278), .ip2(\cache_data_B[7][35] ), .ip3(
        n10172), .ip4(n10171), .op(n10174) );
  nand2_1 U12969 ( .ip1(n11304), .ip2(\cache_data_B[5][35] ), .op(n10173) );
  nand3_1 U12970 ( .ip1(n10175), .ip2(n10174), .ip3(n10173), .op(n12669) );
  nand2_1 U12971 ( .ip1(n12563), .ip2(n12669), .op(n10196) );
  nand2_1 U12972 ( .ip1(\cache_data_B[2][99] ), .ip2(n12486), .op(n10184) );
  and2_1 U12973 ( .ip1(n12582), .ip2(\cache_data_B[5][99] ), .op(n10181) );
  nand2_1 U12974 ( .ip1(n11071), .ip2(\cache_data_B[0][99] ), .op(n10179) );
  nand2_1 U12975 ( .ip1(n12096), .ip2(\cache_data_B[3][99] ), .op(n10178) );
  nand2_1 U12976 ( .ip1(n12371), .ip2(\cache_data_B[6][99] ), .op(n10177) );
  nand2_1 U12977 ( .ip1(n11724), .ip2(\cache_data_B[1][99] ), .op(n10176) );
  nand4_1 U12978 ( .ip1(n10179), .ip2(n10178), .ip3(n10177), .ip4(n10176), 
        .op(n10180) );
  not_ab_or_c_or_d U12979 ( .ip1(\cache_data_B[7][99] ), .ip2(n10575), .ip3(
        n10181), .ip4(n10180), .op(n10183) );
  nand2_1 U12980 ( .ip1(n12054), .ip2(\cache_data_B[4][99] ), .op(n10182) );
  nand3_1 U12981 ( .ip1(n10184), .ip2(n10183), .ip3(n10182), .op(n12658) );
  nand2_1 U12982 ( .ip1(n12573), .ip2(n12658), .op(n10195) );
  nand2_1 U12983 ( .ip1(n10426), .ip2(\cache_data_A[2][99] ), .op(n10193) );
  and2_1 U12984 ( .ip1(n12371), .ip2(\cache_data_A[6][99] ), .op(n10190) );
  nand2_1 U12985 ( .ip1(n12054), .ip2(\cache_data_A[4][99] ), .op(n10188) );
  nand2_1 U12986 ( .ip1(n12096), .ip2(\cache_data_A[3][99] ), .op(n10187) );
  nand2_1 U12987 ( .ip1(n11724), .ip2(\cache_data_A[1][99] ), .op(n10186) );
  nand2_1 U12988 ( .ip1(n11071), .ip2(\cache_data_A[0][99] ), .op(n10185) );
  nand4_1 U12989 ( .ip1(n10188), .ip2(n10187), .ip3(n10186), .ip4(n10185), 
        .op(n10189) );
  not_ab_or_c_or_d U12990 ( .ip1(\cache_data_A[7][99] ), .ip2(n10575), .ip3(
        n10190), .ip4(n10189), .op(n10192) );
  nand2_1 U12991 ( .ip1(n11280), .ip2(\cache_data_A[5][99] ), .op(n10191) );
  nand3_1 U12992 ( .ip1(n10193), .ip2(n10192), .ip3(n10191), .op(n12656) );
  nand2_1 U12993 ( .ip1(n12509), .ip2(n12656), .op(n10194) );
  nand4_1 U12994 ( .ip1(n10197), .ip2(n10196), .ip3(n10195), .ip4(n10194), 
        .op(n10198) );
  not_ab_or_c_or_d U12995 ( .ip1(n12539), .ip2(n12659), .ip3(n10199), .ip4(
        n10198), .op(n10210) );
  nand2_1 U12996 ( .ip1(n10575), .ip2(\cache_data_A[7][35] ), .op(n10208) );
  and2_1 U12997 ( .ip1(n12147), .ip2(\cache_data_A[1][35] ), .op(n10205) );
  nand2_1 U12998 ( .ip1(n11071), .ip2(\cache_data_A[0][35] ), .op(n10203) );
  nand2_1 U12999 ( .ip1(n12337), .ip2(\cache_data_A[6][35] ), .op(n10202) );
  nand2_1 U13000 ( .ip1(n12096), .ip2(\cache_data_A[3][35] ), .op(n10201) );
  nand2_1 U13001 ( .ip1(n10426), .ip2(\cache_data_A[2][35] ), .op(n10200) );
  nand4_1 U13002 ( .ip1(n10203), .ip2(n10202), .ip3(n10201), .ip4(n10200), 
        .op(n10204) );
  not_ab_or_c_or_d U13003 ( .ip1(\cache_data_A[4][35] ), .ip2(n11324), .ip3(
        n10205), .ip4(n10204), .op(n10207) );
  nand2_1 U13004 ( .ip1(n11296), .ip2(\cache_data_A[5][35] ), .op(n10206) );
  nand3_1 U13005 ( .ip1(n10208), .ip2(n10207), .ip3(n10206), .op(n12660) );
  nand2_1 U13006 ( .ip1(n12595), .ip2(n12660), .op(n10209) );
  nand3_1 U13007 ( .ip1(n10211), .ip2(n10210), .ip3(n10209), .op(n10212) );
  mux2_1 U13008 ( .ip1(N4195), .ip2(n10212), .s(n10378), .op(n5317) );
  nand2_1 U13009 ( .ip1(n10426), .ip2(\cache_data_A[2][100] ), .op(n10221) );
  and2_1 U13010 ( .ip1(n11946), .ip2(\cache_data_A[1][100] ), .op(n10218) );
  nand2_1 U13011 ( .ip1(n11296), .ip2(\cache_data_A[5][100] ), .op(n10216) );
  nand2_1 U13012 ( .ip1(n12054), .ip2(\cache_data_A[4][100] ), .op(n10215) );
  nand2_1 U13013 ( .ip1(n12096), .ip2(\cache_data_A[3][100] ), .op(n10214) );
  nand2_1 U13014 ( .ip1(n11071), .ip2(\cache_data_A[0][100] ), .op(n10213) );
  nand4_1 U13015 ( .ip1(n10216), .ip2(n10215), .ip3(n10214), .ip4(n10213), 
        .op(n10217) );
  not_ab_or_c_or_d U13016 ( .ip1(\cache_data_A[7][100] ), .ip2(n10702), .ip3(
        n10218), .ip4(n10217), .op(n10220) );
  nand2_1 U13017 ( .ip1(n12337), .ip2(\cache_data_A[6][100] ), .op(n10219) );
  nand3_1 U13018 ( .ip1(n10221), .ip2(n10220), .ip3(n10219), .op(n12677) );
  nand2_1 U13019 ( .ip1(n12509), .ip2(n12677), .op(n10294) );
  nand2_1 U13020 ( .ip1(n12337), .ip2(\cache_data_A[6][4] ), .op(n10230) );
  and2_1 U13021 ( .ip1(n12410), .ip2(\cache_data_A[3][4] ), .op(n10227) );
  nand2_1 U13022 ( .ip1(n10702), .ip2(\cache_data_A[7][4] ), .op(n10225) );
  nand2_1 U13023 ( .ip1(n10426), .ip2(\cache_data_A[2][4] ), .op(n10224) );
  nand2_1 U13024 ( .ip1(n11304), .ip2(\cache_data_A[5][4] ), .op(n10223) );
  nand2_1 U13025 ( .ip1(n12054), .ip2(\cache_data_A[4][4] ), .op(n10222) );
  nand4_1 U13026 ( .ip1(n10225), .ip2(n10224), .ip3(n10223), .ip4(n10222), 
        .op(n10226) );
  not_ab_or_c_or_d U13027 ( .ip1(\cache_data_A[0][4] ), .ip2(n8452), .ip3(
        n10227), .ip4(n10226), .op(n10229) );
  nand2_1 U13028 ( .ip1(n11724), .ip2(\cache_data_A[1][4] ), .op(n10228) );
  nand3_1 U13029 ( .ip1(n10230), .ip2(n10229), .ip3(n10228), .op(n12674) );
  nand2_1 U13030 ( .ip1(n11057), .ip2(\cache_data_A[7][68] ), .op(n10234) );
  nand2_1 U13031 ( .ip1(n12559), .ip2(\cache_data_A[3][68] ), .op(n10233) );
  nand2_1 U13032 ( .ip1(n12054), .ip2(\cache_data_A[4][68] ), .op(n10232) );
  nand2_1 U13033 ( .ip1(n11724), .ip2(\cache_data_A[1][68] ), .op(n10231) );
  nand4_1 U13034 ( .ip1(n10234), .ip2(n10233), .ip3(n10232), .ip4(n10231), 
        .op(n10240) );
  nand2_1 U13035 ( .ip1(n12337), .ip2(\cache_data_A[6][68] ), .op(n10238) );
  nand2_1 U13036 ( .ip1(n10426), .ip2(\cache_data_A[2][68] ), .op(n10237) );
  nand2_1 U13037 ( .ip1(n11071), .ip2(\cache_data_A[0][68] ), .op(n10236) );
  nand2_1 U13038 ( .ip1(n11304), .ip2(\cache_data_A[5][68] ), .op(n10235) );
  nand4_1 U13039 ( .ip1(n10238), .ip2(n10237), .ip3(n10236), .ip4(n10235), 
        .op(n10239) );
  nor2_1 U13040 ( .ip1(n10240), .ip2(n10239), .op(n12675) );
  nor2_1 U13041 ( .ip1(n12675), .ip2(n12529), .op(n10282) );
  nand2_1 U13042 ( .ip1(n11071), .ip2(\cache_data_B[0][4] ), .op(n10249) );
  and2_1 U13043 ( .ip1(n12476), .ip2(\cache_data_B[4][4] ), .op(n10246) );
  nand2_1 U13044 ( .ip1(n10686), .ip2(\cache_data_B[1][4] ), .op(n10244) );
  nand2_1 U13045 ( .ip1(n12337), .ip2(\cache_data_B[6][4] ), .op(n10243) );
  nand2_1 U13046 ( .ip1(n12096), .ip2(\cache_data_B[3][4] ), .op(n10242) );
  nand2_1 U13047 ( .ip1(n10702), .ip2(\cache_data_B[7][4] ), .op(n10241) );
  nand4_1 U13048 ( .ip1(n10244), .ip2(n10243), .ip3(n10242), .ip4(n10241), 
        .op(n10245) );
  not_ab_or_c_or_d U13049 ( .ip1(\cache_data_B[2][4] ), .ip2(n12546), .ip3(
        n10246), .ip4(n10245), .op(n10248) );
  nand2_1 U13050 ( .ip1(n11280), .ip2(\cache_data_B[5][4] ), .op(n10247) );
  nand3_1 U13051 ( .ip1(n10249), .ip2(n10248), .ip3(n10247), .op(n12679) );
  nand2_1 U13052 ( .ip1(n12539), .ip2(n12679), .op(n10280) );
  nand2_1 U13053 ( .ip1(n12337), .ip2(\cache_data_B[6][36] ), .op(n10258) );
  and2_1 U13054 ( .ip1(n12581), .ip2(\cache_data_B[7][36] ), .op(n10255) );
  nand2_1 U13055 ( .ip1(n11236), .ip2(\cache_data_B[5][36] ), .op(n10253) );
  nand2_1 U13056 ( .ip1(n10426), .ip2(\cache_data_B[2][36] ), .op(n10252) );
  nand2_1 U13057 ( .ip1(n10686), .ip2(\cache_data_B[1][36] ), .op(n10251) );
  nand2_1 U13058 ( .ip1(n12096), .ip2(\cache_data_B[3][36] ), .op(n10250) );
  nand4_1 U13059 ( .ip1(n10253), .ip2(n10252), .ip3(n10251), .ip4(n10250), 
        .op(n10254) );
  not_ab_or_c_or_d U13060 ( .ip1(\cache_data_B[0][36] ), .ip2(n11911), .ip3(
        n10255), .ip4(n10254), .op(n10257) );
  nand2_1 U13061 ( .ip1(n11324), .ip2(\cache_data_B[4][36] ), .op(n10256) );
  nand3_1 U13062 ( .ip1(n10258), .ip2(n10257), .ip3(n10256), .op(n12678) );
  nand2_1 U13063 ( .ip1(n12563), .ip2(n12678), .op(n10279) );
  nand2_1 U13064 ( .ip1(\cache_data_B[6][100] ), .ip2(n12371), .op(n10267) );
  and2_1 U13065 ( .ip1(n8060), .ip2(\cache_data_B[3][100] ), .op(n10264) );
  nand2_1 U13066 ( .ip1(n10686), .ip2(\cache_data_B[1][100] ), .op(n10262) );
  nand2_1 U13067 ( .ip1(n11071), .ip2(\cache_data_B[0][100] ), .op(n10261) );
  nand2_1 U13068 ( .ip1(n10575), .ip2(\cache_data_B[7][100] ), .op(n10260) );
  nand2_1 U13069 ( .ip1(n11236), .ip2(\cache_data_B[5][100] ), .op(n10259) );
  nand4_1 U13070 ( .ip1(n10262), .ip2(n10261), .ip3(n10260), .ip4(n10259), 
        .op(n10263) );
  not_ab_or_c_or_d U13071 ( .ip1(n12546), .ip2(\cache_data_B[2][100] ), .ip3(
        n10264), .ip4(n10263), .op(n10266) );
  nand2_1 U13072 ( .ip1(n11324), .ip2(\cache_data_B[4][100] ), .op(n10265) );
  nand3_1 U13073 ( .ip1(n10267), .ip2(n10266), .ip3(n10265), .op(n12676) );
  nand2_1 U13074 ( .ip1(n12573), .ip2(n12676), .op(n10278) );
  nand2_1 U13075 ( .ip1(n10426), .ip2(\cache_data_B[2][68] ), .op(n10276) );
  and2_1 U13076 ( .ip1(n11156), .ip2(\cache_data_B[4][68] ), .op(n10273) );
  nand2_1 U13077 ( .ip1(n12581), .ip2(\cache_data_B[7][68] ), .op(n10271) );
  nand2_1 U13078 ( .ip1(n12337), .ip2(\cache_data_B[6][68] ), .op(n10270) );
  nand2_1 U13079 ( .ip1(n11296), .ip2(\cache_data_B[5][68] ), .op(n10269) );
  nand2_1 U13080 ( .ip1(n12096), .ip2(\cache_data_B[3][68] ), .op(n10268) );
  nand4_1 U13081 ( .ip1(n10271), .ip2(n10270), .ip3(n10269), .ip4(n10268), 
        .op(n10272) );
  not_ab_or_c_or_d U13082 ( .ip1(n12297), .ip2(\cache_data_B[0][68] ), .ip3(
        n10273), .ip4(n10272), .op(n10275) );
  nand2_1 U13083 ( .ip1(n11724), .ip2(\cache_data_B[1][68] ), .op(n10274) );
  nand3_1 U13084 ( .ip1(n10276), .ip2(n10275), .ip3(n10274), .op(n12686) );
  nand2_1 U13085 ( .ip1(n12580), .ip2(n12686), .op(n10277) );
  nand4_1 U13086 ( .ip1(n10280), .ip2(n10279), .ip3(n10278), .ip4(n10277), 
        .op(n10281) );
  not_ab_or_c_or_d U13087 ( .ip1(n12550), .ip2(n12674), .ip3(n10282), .ip4(
        n10281), .op(n10293) );
  nand2_1 U13088 ( .ip1(\cache_data_A[3][36] ), .ip2(n12410), .op(n10291) );
  and2_1 U13089 ( .ip1(n10166), .ip2(\cache_data_A[1][36] ), .op(n10288) );
  nand2_1 U13090 ( .ip1(n12278), .ip2(\cache_data_A[7][36] ), .op(n10286) );
  nand2_1 U13091 ( .ip1(n11156), .ip2(\cache_data_A[4][36] ), .op(n10285) );
  nand2_1 U13092 ( .ip1(n10426), .ip2(\cache_data_A[2][36] ), .op(n10284) );
  nand2_1 U13093 ( .ip1(n12337), .ip2(\cache_data_A[6][36] ), .op(n10283) );
  nand4_1 U13094 ( .ip1(n10286), .ip2(n10285), .ip3(n10284), .ip4(n10283), 
        .op(n10287) );
  not_ab_or_c_or_d U13095 ( .ip1(n12297), .ip2(\cache_data_A[0][36] ), .ip3(
        n10288), .ip4(n10287), .op(n10290) );
  nand2_1 U13096 ( .ip1(n11236), .ip2(\cache_data_A[5][36] ), .op(n10289) );
  nand3_1 U13097 ( .ip1(n10291), .ip2(n10290), .ip3(n10289), .op(n12687) );
  nand2_1 U13098 ( .ip1(n12595), .ip2(n12687), .op(n10292) );
  nand3_1 U13099 ( .ip1(n10294), .ip2(n10293), .ip3(n10292), .op(n10295) );
  mux2_1 U13100 ( .ip1(N4192), .ip2(n10295), .s(n10378), .op(n5316) );
  nand2_1 U13101 ( .ip1(n12337), .ip2(\cache_data_B[6][101] ), .op(n10304) );
  and2_1 U13102 ( .ip1(n12256), .ip2(\cache_data_B[5][101] ), .op(n10301) );
  nand2_1 U13103 ( .ip1(n10426), .ip2(\cache_data_B[2][101] ), .op(n10299) );
  nand2_1 U13104 ( .ip1(n12278), .ip2(\cache_data_B[7][101] ), .op(n10298) );
  nand2_1 U13105 ( .ip1(n11071), .ip2(\cache_data_B[0][101] ), .op(n10297) );
  nand2_1 U13106 ( .ip1(n10686), .ip2(\cache_data_B[1][101] ), .op(n10296) );
  nand4_1 U13107 ( .ip1(n10299), .ip2(n10298), .ip3(n10297), .ip4(n10296), 
        .op(n10300) );
  not_ab_or_c_or_d U13108 ( .ip1(n11156), .ip2(\cache_data_B[4][101] ), .ip3(
        n10301), .ip4(n10300), .op(n10303) );
  nand2_1 U13109 ( .ip1(n12559), .ip2(\cache_data_B[3][101] ), .op(n10302) );
  nand3_1 U13110 ( .ip1(n10304), .ip2(n10303), .ip3(n10302), .op(n12694) );
  nand2_1 U13111 ( .ip1(n12573), .ip2(n12694), .op(n10377) );
  nand2_1 U13112 ( .ip1(n12337), .ip2(\cache_data_A[6][5] ), .op(n10313) );
  and2_1 U13113 ( .ip1(n12468), .ip2(\cache_data_A[7][5] ), .op(n10310) );
  nand2_1 U13114 ( .ip1(n10686), .ip2(\cache_data_A[1][5] ), .op(n10308) );
  nand2_1 U13115 ( .ip1(n12559), .ip2(\cache_data_A[3][5] ), .op(n10307) );
  nand2_1 U13116 ( .ip1(n11296), .ip2(\cache_data_A[5][5] ), .op(n10306) );
  nand2_1 U13117 ( .ip1(n10426), .ip2(\cache_data_A[2][5] ), .op(n10305) );
  nand4_1 U13118 ( .ip1(n10308), .ip2(n10307), .ip3(n10306), .ip4(n10305), 
        .op(n10309) );
  not_ab_or_c_or_d U13119 ( .ip1(n12297), .ip2(\cache_data_A[0][5] ), .ip3(
        n10310), .ip4(n10309), .op(n10312) );
  nand2_1 U13120 ( .ip1(n11156), .ip2(\cache_data_A[4][5] ), .op(n10311) );
  nand3_1 U13121 ( .ip1(n10313), .ip2(n10312), .ip3(n10311), .op(n12692) );
  nand2_1 U13122 ( .ip1(n12559), .ip2(\cache_data_A[3][69] ), .op(n10317) );
  nand2_1 U13123 ( .ip1(n12278), .ip2(\cache_data_A[7][69] ), .op(n10316) );
  nand2_1 U13124 ( .ip1(n11324), .ip2(\cache_data_A[4][69] ), .op(n10315) );
  nand2_1 U13125 ( .ip1(n11724), .ip2(\cache_data_A[1][69] ), .op(n10314) );
  nand4_1 U13126 ( .ip1(n10317), .ip2(n10316), .ip3(n10315), .ip4(n10314), 
        .op(n10323) );
  nand2_1 U13127 ( .ip1(n11071), .ip2(\cache_data_A[0][69] ), .op(n10321) );
  nand2_1 U13128 ( .ip1(n12337), .ip2(\cache_data_A[6][69] ), .op(n10320) );
  nand2_1 U13129 ( .ip1(n11280), .ip2(\cache_data_A[5][69] ), .op(n10319) );
  nand2_1 U13130 ( .ip1(n10426), .ip2(\cache_data_A[2][69] ), .op(n10318) );
  nand4_1 U13131 ( .ip1(n10321), .ip2(n10320), .ip3(n10319), .ip4(n10318), 
        .op(n10322) );
  nor2_1 U13132 ( .ip1(n10323), .ip2(n10322), .op(n12693) );
  nor2_1 U13133 ( .ip1(n12693), .ip2(n12529), .op(n10365) );
  nand2_1 U13134 ( .ip1(n12559), .ip2(\cache_data_A[3][101] ), .op(n10332) );
  and2_1 U13135 ( .ip1(n11296), .ip2(\cache_data_A[5][101] ), .op(n10329) );
  nand2_1 U13136 ( .ip1(n10426), .ip2(\cache_data_A[2][101] ), .op(n10327) );
  nand2_1 U13137 ( .ip1(n12278), .ip2(\cache_data_A[7][101] ), .op(n10326) );
  nand2_1 U13138 ( .ip1(n11324), .ip2(\cache_data_A[4][101] ), .op(n10325) );
  nand2_1 U13139 ( .ip1(n11071), .ip2(\cache_data_A[0][101] ), .op(n10324) );
  nand4_1 U13140 ( .ip1(n10327), .ip2(n10326), .ip3(n10325), .ip4(n10324), 
        .op(n10328) );
  not_ab_or_c_or_d U13141 ( .ip1(\cache_data_A[6][101] ), .ip2(n12551), .ip3(
        n10329), .ip4(n10328), .op(n10331) );
  nand2_1 U13142 ( .ip1(n11724), .ip2(\cache_data_A[1][101] ), .op(n10330) );
  nand3_1 U13143 ( .ip1(n10332), .ip2(n10331), .ip3(n10330), .op(n12704) );
  nand2_1 U13144 ( .ip1(n12509), .ip2(n12704), .op(n10363) );
  nand2_1 U13145 ( .ip1(\cache_data_B[4][37] ), .ip2(n12194), .op(n10341) );
  and2_1 U13146 ( .ip1(n12582), .ip2(\cache_data_B[5][37] ), .op(n10338) );
  nand2_1 U13147 ( .ip1(n10575), .ip2(\cache_data_B[7][37] ), .op(n10336) );
  nand2_1 U13148 ( .ip1(n12096), .ip2(\cache_data_B[3][37] ), .op(n10335) );
  nand2_1 U13149 ( .ip1(n10426), .ip2(\cache_data_B[2][37] ), .op(n10334) );
  nand2_1 U13150 ( .ip1(n12337), .ip2(\cache_data_B[6][37] ), .op(n10333) );
  nand4_1 U13151 ( .ip1(n10336), .ip2(n10335), .ip3(n10334), .ip4(n10333), 
        .op(n10337) );
  not_ab_or_c_or_d U13152 ( .ip1(n12204), .ip2(\cache_data_B[0][37] ), .ip3(
        n10338), .ip4(n10337), .op(n10340) );
  nand2_1 U13153 ( .ip1(n10686), .ip2(\cache_data_B[1][37] ), .op(n10339) );
  nand3_1 U13154 ( .ip1(n10341), .ip2(n10340), .ip3(n10339), .op(n12697) );
  nand2_1 U13155 ( .ip1(n12563), .ip2(n12697), .op(n10362) );
  nand2_1 U13156 ( .ip1(n12278), .ip2(\cache_data_B[7][5] ), .op(n10350) );
  and2_1 U13157 ( .ip1(n12582), .ip2(\cache_data_B[5][5] ), .op(n10347) );
  nand2_1 U13158 ( .ip1(n11535), .ip2(\cache_data_B[3][5] ), .op(n10345) );
  nand2_1 U13159 ( .ip1(n10686), .ip2(\cache_data_B[1][5] ), .op(n10344) );
  nand2_1 U13160 ( .ip1(n11071), .ip2(\cache_data_B[0][5] ), .op(n10343) );
  nand2_1 U13161 ( .ip1(n10426), .ip2(\cache_data_B[2][5] ), .op(n10342) );
  nand4_1 U13162 ( .ip1(n10345), .ip2(n10344), .ip3(n10343), .ip4(n10342), 
        .op(n10346) );
  not_ab_or_c_or_d U13163 ( .ip1(n12551), .ip2(\cache_data_B[6][5] ), .ip3(
        n10347), .ip4(n10346), .op(n10349) );
  nand2_1 U13164 ( .ip1(n12054), .ip2(\cache_data_B[4][5] ), .op(n10348) );
  nand3_1 U13165 ( .ip1(n10350), .ip2(n10349), .ip3(n10348), .op(n12695) );
  nand2_1 U13166 ( .ip1(n12539), .ip2(n12695), .op(n10361) );
  nand2_1 U13167 ( .ip1(n12559), .ip2(\cache_data_A[3][37] ), .op(n10359) );
  and2_1 U13168 ( .ip1(n12458), .ip2(\cache_data_A[6][37] ), .op(n10356) );
  nand2_1 U13169 ( .ip1(n10686), .ip2(\cache_data_A[1][37] ), .op(n10354) );
  nand2_1 U13170 ( .ip1(n10426), .ip2(\cache_data_A[2][37] ), .op(n10353) );
  nand2_1 U13171 ( .ip1(n11071), .ip2(\cache_data_A[0][37] ), .op(n10352) );
  nand2_1 U13172 ( .ip1(n11236), .ip2(\cache_data_A[5][37] ), .op(n10351) );
  nand4_1 U13173 ( .ip1(n10354), .ip2(n10353), .ip3(n10352), .ip4(n10351), 
        .op(n10355) );
  not_ab_or_c_or_d U13174 ( .ip1(n12552), .ip2(\cache_data_A[7][37] ), .ip3(
        n10356), .ip4(n10355), .op(n10358) );
  nand2_1 U13175 ( .ip1(n11156), .ip2(\cache_data_A[4][37] ), .op(n10357) );
  nand3_1 U13176 ( .ip1(n10359), .ip2(n10358), .ip3(n10357), .op(n12705) );
  nand2_1 U13177 ( .ip1(n12595), .ip2(n12705), .op(n10360) );
  nand4_1 U13178 ( .ip1(n10363), .ip2(n10362), .ip3(n10361), .ip4(n10360), 
        .op(n10364) );
  not_ab_or_c_or_d U13179 ( .ip1(n12550), .ip2(n12692), .ip3(n10365), .ip4(
        n10364), .op(n10376) );
  nand2_1 U13180 ( .ip1(n10426), .ip2(\cache_data_B[2][69] ), .op(n10374) );
  and2_1 U13181 ( .ip1(n11156), .ip2(\cache_data_B[4][69] ), .op(n10371) );
  nand2_1 U13182 ( .ip1(n12278), .ip2(\cache_data_B[7][69] ), .op(n10369) );
  nand2_1 U13183 ( .ip1(n11071), .ip2(\cache_data_B[0][69] ), .op(n10368) );
  nand2_1 U13184 ( .ip1(n11236), .ip2(\cache_data_B[5][69] ), .op(n10367) );
  nand2_1 U13185 ( .ip1(n10686), .ip2(\cache_data_B[1][69] ), .op(n10366) );
  nand4_1 U13186 ( .ip1(n10369), .ip2(n10368), .ip3(n10367), .ip4(n10366), 
        .op(n10370) );
  not_ab_or_c_or_d U13187 ( .ip1(\cache_data_B[3][69] ), .ip2(n11535), .ip3(
        n10371), .ip4(n10370), .op(n10373) );
  nand2_1 U13188 ( .ip1(n12337), .ip2(\cache_data_B[6][69] ), .op(n10372) );
  nand3_1 U13189 ( .ip1(n10374), .ip2(n10373), .ip3(n10372), .op(n12696) );
  nand2_1 U13190 ( .ip1(n12580), .ip2(n12696), .op(n10375) );
  nand3_1 U13191 ( .ip1(n10377), .ip2(n10376), .ip3(n10375), .op(n10379) );
  mux2_1 U13192 ( .ip1(N4189), .ip2(n10379), .s(n10378), .op(n5315) );
  nand2_1 U13193 ( .ip1(n11071), .ip2(\cache_data_B[0][102] ), .op(n10388) );
  and2_1 U13194 ( .ip1(n11296), .ip2(\cache_data_B[5][102] ), .op(n10385) );
  nand2_1 U13195 ( .ip1(n12337), .ip2(\cache_data_B[6][102] ), .op(n10383) );
  nand2_1 U13196 ( .ip1(n12054), .ip2(\cache_data_B[4][102] ), .op(n10382) );
  nand2_1 U13197 ( .ip1(n11535), .ip2(\cache_data_B[3][102] ), .op(n10381) );
  nand2_1 U13198 ( .ip1(n10575), .ip2(\cache_data_B[7][102] ), .op(n10380) );
  nand4_1 U13199 ( .ip1(n10383), .ip2(n10382), .ip3(n10381), .ip4(n10380), 
        .op(n10384) );
  not_ab_or_c_or_d U13200 ( .ip1(\cache_data_B[2][102] ), .ip2(n12546), .ip3(
        n10385), .ip4(n10384), .op(n10387) );
  nand2_1 U13201 ( .ip1(n11724), .ip2(\cache_data_B[1][102] ), .op(n10386) );
  nand3_1 U13202 ( .ip1(n10388), .ip2(n10387), .ip3(n10386), .op(n12712) );
  nand2_1 U13203 ( .ip1(n12573), .ip2(n12712), .op(n10462) );
  nand2_1 U13204 ( .ip1(\cache_data_B[0][38] ), .ip2(n12370), .op(n10397) );
  and2_1 U13205 ( .ip1(n12147), .ip2(\cache_data_B[1][38] ), .op(n10394) );
  nand2_1 U13206 ( .ip1(n11535), .ip2(\cache_data_B[3][38] ), .op(n10392) );
  nand2_1 U13207 ( .ip1(n11236), .ip2(\cache_data_B[5][38] ), .op(n10391) );
  nand2_1 U13208 ( .ip1(n12278), .ip2(\cache_data_B[7][38] ), .op(n10390) );
  nand2_1 U13209 ( .ip1(n12320), .ip2(\cache_data_B[6][38] ), .op(n10389) );
  nand4_1 U13210 ( .ip1(n10392), .ip2(n10391), .ip3(n10390), .ip4(n10389), 
        .op(n10393) );
  not_ab_or_c_or_d U13211 ( .ip1(n12546), .ip2(\cache_data_B[2][38] ), .ip3(
        n10394), .ip4(n10393), .op(n10396) );
  nand2_1 U13212 ( .ip1(n11324), .ip2(\cache_data_B[4][38] ), .op(n10395) );
  nand3_1 U13213 ( .ip1(n10397), .ip2(n10396), .ip3(n10395), .op(n12715) );
  nand2_1 U13214 ( .ip1(n12278), .ip2(\cache_data_A[7][70] ), .op(n10401) );
  nand2_1 U13215 ( .ip1(n11071), .ip2(\cache_data_A[0][70] ), .op(n10400) );
  nand2_1 U13216 ( .ip1(n10426), .ip2(\cache_data_A[2][70] ), .op(n10399) );
  nand2_1 U13217 ( .ip1(n11296), .ip2(\cache_data_A[5][70] ), .op(n10398) );
  nand4_1 U13218 ( .ip1(n10401), .ip2(n10400), .ip3(n10399), .ip4(n10398), 
        .op(n10407) );
  nand2_1 U13219 ( .ip1(n12559), .ip2(\cache_data_A[3][70] ), .op(n10405) );
  nand2_1 U13220 ( .ip1(n12371), .ip2(\cache_data_A[6][70] ), .op(n10404) );
  nand2_1 U13221 ( .ip1(n11156), .ip2(\cache_data_A[4][70] ), .op(n10403) );
  nand2_1 U13222 ( .ip1(n11724), .ip2(\cache_data_A[1][70] ), .op(n10402) );
  nand4_1 U13223 ( .ip1(n10405), .ip2(n10404), .ip3(n10403), .ip4(n10402), 
        .op(n10406) );
  nor2_1 U13224 ( .ip1(n10407), .ip2(n10406), .op(n12711) );
  nor2_1 U13225 ( .ip1(n12711), .ip2(n12529), .op(n10450) );
  nand2_1 U13226 ( .ip1(n12320), .ip2(\cache_data_A[6][102] ), .op(n10416) );
  and2_1 U13227 ( .ip1(n12582), .ip2(\cache_data_A[5][102] ), .op(n10413) );
  nand2_1 U13228 ( .ip1(n11724), .ip2(\cache_data_A[1][102] ), .op(n10411) );
  nand2_1 U13229 ( .ip1(n12054), .ip2(\cache_data_A[4][102] ), .op(n10410) );
  nand2_1 U13230 ( .ip1(n10426), .ip2(\cache_data_A[2][102] ), .op(n10409) );
  nand2_1 U13231 ( .ip1(n10575), .ip2(\cache_data_A[7][102] ), .op(n10408) );
  nand4_1 U13232 ( .ip1(n10411), .ip2(n10410), .ip3(n10409), .ip4(n10408), 
        .op(n10412) );
  not_ab_or_c_or_d U13233 ( .ip1(n12297), .ip2(\cache_data_A[0][102] ), .ip3(
        n10413), .ip4(n10412), .op(n10415) );
  nand2_1 U13234 ( .ip1(n12559), .ip2(\cache_data_A[3][102] ), .op(n10414) );
  nand3_1 U13235 ( .ip1(n10416), .ip2(n10415), .ip3(n10414), .op(n12714) );
  nand2_1 U13236 ( .ip1(n12509), .ip2(n12714), .op(n10448) );
  nand2_1 U13237 ( .ip1(n12278), .ip2(\cache_data_B[7][6] ), .op(n10425) );
  and2_1 U13238 ( .ip1(n12582), .ip2(\cache_data_B[5][6] ), .op(n10422) );
  nand2_1 U13239 ( .ip1(n12559), .ip2(\cache_data_B[3][6] ), .op(n10420) );
  nand2_1 U13240 ( .ip1(n11724), .ip2(\cache_data_B[1][6] ), .op(n10419) );
  nand2_1 U13241 ( .ip1(n11071), .ip2(\cache_data_B[0][6] ), .op(n10418) );
  nand2_1 U13242 ( .ip1(n10426), .ip2(\cache_data_B[2][6] ), .op(n10417) );
  nand4_1 U13243 ( .ip1(n10420), .ip2(n10419), .ip3(n10418), .ip4(n10417), 
        .op(n10421) );
  not_ab_or_c_or_d U13244 ( .ip1(\cache_data_B[4][6] ), .ip2(n11156), .ip3(
        n10422), .ip4(n10421), .op(n10424) );
  nand2_1 U13245 ( .ip1(n12458), .ip2(\cache_data_B[6][6] ), .op(n10423) );
  nand3_1 U13246 ( .ip1(n10425), .ip2(n10424), .ip3(n10423), .op(n12722) );
  nand2_1 U13247 ( .ip1(n12539), .ip2(n12722), .op(n10447) );
  nand2_1 U13248 ( .ip1(n10426), .ip2(\cache_data_B[2][70] ), .op(n10435) );
  and2_1 U13249 ( .ip1(n12582), .ip2(\cache_data_B[5][70] ), .op(n10432) );
  nand2_1 U13250 ( .ip1(n12320), .ip2(\cache_data_B[6][70] ), .op(n10430) );
  nand2_1 U13251 ( .ip1(n10575), .ip2(\cache_data_B[7][70] ), .op(n10429) );
  nand2_1 U13252 ( .ip1(n10686), .ip2(\cache_data_B[1][70] ), .op(n10428) );
  nand2_1 U13253 ( .ip1(n12584), .ip2(\cache_data_B[4][70] ), .op(n10427) );
  nand4_1 U13254 ( .ip1(n10430), .ip2(n10429), .ip3(n10428), .ip4(n10427), 
        .op(n10431) );
  not_ab_or_c_or_d U13255 ( .ip1(\cache_data_B[0][70] ), .ip2(n11911), .ip3(
        n10432), .ip4(n10431), .op(n10434) );
  nand2_1 U13256 ( .ip1(n11535), .ip2(\cache_data_B[3][70] ), .op(n10433) );
  nand3_1 U13257 ( .ip1(n10435), .ip2(n10434), .ip3(n10433), .op(n12713) );
  nand2_1 U13258 ( .ip1(n12580), .ip2(n12713), .op(n10446) );
  nand2_1 U13259 ( .ip1(\cache_data_A[7][6] ), .ip2(n12552), .op(n10444) );
  and2_1 U13260 ( .ip1(n12147), .ip2(\cache_data_A[1][6] ), .op(n10441) );
  nand2_1 U13261 ( .ip1(n11142), .ip2(\cache_data_A[2][6] ), .op(n10439) );
  nand2_1 U13262 ( .ip1(n11071), .ip2(\cache_data_A[0][6] ), .op(n10438) );
  nand2_1 U13263 ( .ip1(n11780), .ip2(\cache_data_A[6][6] ), .op(n10437) );
  nand2_1 U13264 ( .ip1(n12584), .ip2(\cache_data_A[4][6] ), .op(n10436) );
  nand4_1 U13265 ( .ip1(n10439), .ip2(n10438), .ip3(n10437), .ip4(n10436), 
        .op(n10440) );
  not_ab_or_c_or_d U13266 ( .ip1(\cache_data_A[3][6] ), .ip2(n12559), .ip3(
        n10441), .ip4(n10440), .op(n10443) );
  nand2_1 U13267 ( .ip1(n11296), .ip2(\cache_data_A[5][6] ), .op(n10442) );
  nand3_1 U13268 ( .ip1(n10444), .ip2(n10443), .ip3(n10442), .op(n12710) );
  nand2_1 U13269 ( .ip1(n12550), .ip2(n12710), .op(n10445) );
  nand4_1 U13270 ( .ip1(n10448), .ip2(n10447), .ip3(n10446), .ip4(n10445), 
        .op(n10449) );
  not_ab_or_c_or_d U13271 ( .ip1(n12563), .ip2(n12715), .ip3(n10450), .ip4(
        n10449), .op(n10461) );
  nand2_1 U13272 ( .ip1(\cache_data_A[3][38] ), .ip2(n12410), .op(n10459) );
  and2_1 U13273 ( .ip1(n12486), .ip2(\cache_data_A[2][38] ), .op(n10456) );
  nand2_1 U13274 ( .ip1(n10575), .ip2(\cache_data_A[7][38] ), .op(n10454) );
  nand2_1 U13275 ( .ip1(n11296), .ip2(\cache_data_A[5][38] ), .op(n10453) );
  nand2_1 U13276 ( .ip1(n11156), .ip2(\cache_data_A[4][38] ), .op(n10452) );
  nand2_1 U13277 ( .ip1(n12458), .ip2(\cache_data_A[6][38] ), .op(n10451) );
  nand4_1 U13278 ( .ip1(n10454), .ip2(n10453), .ip3(n10452), .ip4(n10451), 
        .op(n10455) );
  not_ab_or_c_or_d U13279 ( .ip1(n12297), .ip2(\cache_data_A[0][38] ), .ip3(
        n10456), .ip4(n10455), .op(n10458) );
  nand2_1 U13280 ( .ip1(n11724), .ip2(\cache_data_A[1][38] ), .op(n10457) );
  nand3_1 U13281 ( .ip1(n10459), .ip2(n10458), .ip3(n10457), .op(n12723) );
  nand2_1 U13282 ( .ip1(n12595), .ip2(n12723), .op(n10460) );
  nand3_1 U13283 ( .ip1(n10462), .ip2(n10461), .ip3(n10460), .op(n10463) );
  mux2_1 U13284 ( .ip1(N4186), .ip2(n10463), .s(n11472), .op(n5314) );
  nand2_1 U13285 ( .ip1(n11142), .ip2(\cache_data_A[2][103] ), .op(n10472) );
  and2_1 U13286 ( .ip1(n11156), .ip2(\cache_data_A[4][103] ), .op(n10469) );
  nand2_1 U13287 ( .ip1(n11296), .ip2(\cache_data_A[5][103] ), .op(n10467) );
  nand2_1 U13288 ( .ip1(n11780), .ip2(\cache_data_A[6][103] ), .op(n10466) );
  nand2_1 U13289 ( .ip1(n12559), .ip2(\cache_data_A[3][103] ), .op(n10465) );
  nand2_1 U13290 ( .ip1(n11071), .ip2(\cache_data_A[0][103] ), .op(n10464) );
  nand4_1 U13291 ( .ip1(n10467), .ip2(n10466), .ip3(n10465), .ip4(n10464), 
        .op(n10468) );
  not_ab_or_c_or_d U13292 ( .ip1(n12278), .ip2(\cache_data_A[7][103] ), .ip3(
        n10469), .ip4(n10468), .op(n10471) );
  nand2_1 U13293 ( .ip1(n11724), .ip2(\cache_data_A[1][103] ), .op(n10470) );
  nand3_1 U13294 ( .ip1(n10472), .ip2(n10471), .ip3(n10470), .op(n12740) );
  nand2_1 U13295 ( .ip1(n12509), .ip2(n12740), .op(n10545) );
  nand2_1 U13296 ( .ip1(n10575), .ip2(\cache_data_A[7][7] ), .op(n10481) );
  and2_1 U13297 ( .ip1(n12147), .ip2(\cache_data_A[1][7] ), .op(n10478) );
  nand2_1 U13298 ( .ip1(n12559), .ip2(\cache_data_A[3][7] ), .op(n10476) );
  nand2_1 U13299 ( .ip1(n12054), .ip2(\cache_data_A[4][7] ), .op(n10475) );
  nand2_1 U13300 ( .ip1(n11071), .ip2(\cache_data_A[0][7] ), .op(n10474) );
  nand2_1 U13301 ( .ip1(n11142), .ip2(\cache_data_A[2][7] ), .op(n10473) );
  nand4_1 U13302 ( .ip1(n10476), .ip2(n10475), .ip3(n10474), .ip4(n10473), 
        .op(n10477) );
  not_ab_or_c_or_d U13303 ( .ip1(\cache_data_A[6][7] ), .ip2(n12551), .ip3(
        n10478), .ip4(n10477), .op(n10480) );
  nand2_1 U13304 ( .ip1(n11296), .ip2(\cache_data_A[5][7] ), .op(n10479) );
  nand3_1 U13305 ( .ip1(n10481), .ip2(n10480), .ip3(n10479), .op(n12728) );
  nand2_1 U13306 ( .ip1(n11724), .ip2(\cache_data_A[1][71] ), .op(n10485) );
  nand2_1 U13307 ( .ip1(n12371), .ip2(\cache_data_A[6][71] ), .op(n10484) );
  nand2_1 U13308 ( .ip1(n11142), .ip2(\cache_data_A[2][71] ), .op(n10483) );
  nand2_1 U13309 ( .ip1(n10575), .ip2(\cache_data_A[7][71] ), .op(n10482) );
  nand4_1 U13310 ( .ip1(n10485), .ip2(n10484), .ip3(n10483), .ip4(n10482), 
        .op(n10491) );
  nand2_1 U13311 ( .ip1(n11071), .ip2(\cache_data_A[0][71] ), .op(n10489) );
  nand2_1 U13312 ( .ip1(n12096), .ip2(\cache_data_A[3][71] ), .op(n10488) );
  nand2_1 U13313 ( .ip1(n11296), .ip2(\cache_data_A[5][71] ), .op(n10487) );
  nand2_1 U13314 ( .ip1(n12054), .ip2(\cache_data_A[4][71] ), .op(n10486) );
  nand4_1 U13315 ( .ip1(n10489), .ip2(n10488), .ip3(n10487), .ip4(n10486), 
        .op(n10490) );
  nor2_1 U13316 ( .ip1(n10491), .ip2(n10490), .op(n12729) );
  nor2_1 U13317 ( .ip1(n12729), .ip2(n12529), .op(n10533) );
  nand2_1 U13318 ( .ip1(\cache_data_A[7][39] ), .ip2(n12552), .op(n10500) );
  and2_1 U13319 ( .ip1(n12591), .ip2(\cache_data_A[3][39] ), .op(n10497) );
  nand2_1 U13320 ( .ip1(n12054), .ip2(\cache_data_A[4][39] ), .op(n10495) );
  nand2_1 U13321 ( .ip1(n11142), .ip2(\cache_data_A[2][39] ), .op(n10494) );
  nand2_1 U13322 ( .ip1(n11780), .ip2(\cache_data_A[6][39] ), .op(n10493) );
  nand2_1 U13323 ( .ip1(n10686), .ip2(\cache_data_A[1][39] ), .op(n10492) );
  nand4_1 U13324 ( .ip1(n10495), .ip2(n10494), .ip3(n10493), .ip4(n10492), 
        .op(n10496) );
  not_ab_or_c_or_d U13325 ( .ip1(n12297), .ip2(\cache_data_A[0][39] ), .ip3(
        n10497), .ip4(n10496), .op(n10499) );
  nand2_1 U13326 ( .ip1(n11296), .ip2(\cache_data_A[5][39] ), .op(n10498) );
  nand3_1 U13327 ( .ip1(n10500), .ip2(n10499), .ip3(n10498), .op(n12732) );
  nand2_1 U13328 ( .ip1(n12595), .ip2(n12732), .op(n10531) );
  nand2_1 U13329 ( .ip1(n10575), .ip2(\cache_data_B[7][7] ), .op(n10509) );
  and2_1 U13330 ( .ip1(n12410), .ip2(\cache_data_B[3][7] ), .op(n10506) );
  nand2_1 U13331 ( .ip1(n11236), .ip2(\cache_data_B[5][7] ), .op(n10504) );
  nand2_1 U13332 ( .ip1(n11071), .ip2(\cache_data_B[0][7] ), .op(n10503) );
  nand2_1 U13333 ( .ip1(n12320), .ip2(\cache_data_B[6][7] ), .op(n10502) );
  nand2_1 U13334 ( .ip1(n10686), .ip2(\cache_data_B[1][7] ), .op(n10501) );
  nand4_1 U13335 ( .ip1(n10504), .ip2(n10503), .ip3(n10502), .ip4(n10501), 
        .op(n10505) );
  not_ab_or_c_or_d U13336 ( .ip1(\cache_data_B[2][7] ), .ip2(n12546), .ip3(
        n10506), .ip4(n10505), .op(n10508) );
  nand2_1 U13337 ( .ip1(n12054), .ip2(\cache_data_B[4][7] ), .op(n10507) );
  nand3_1 U13338 ( .ip1(n10509), .ip2(n10508), .ip3(n10507), .op(n12730) );
  nand2_1 U13339 ( .ip1(n12539), .ip2(n12730), .op(n10530) );
  nand2_1 U13340 ( .ip1(n12559), .ip2(\cache_data_B[3][39] ), .op(n10518) );
  and2_1 U13341 ( .ip1(n11296), .ip2(\cache_data_B[5][39] ), .op(n10515) );
  nand2_1 U13342 ( .ip1(n11071), .ip2(\cache_data_B[0][39] ), .op(n10513) );
  nand2_1 U13343 ( .ip1(n10686), .ip2(\cache_data_B[1][39] ), .op(n10512) );
  nand2_1 U13344 ( .ip1(n11142), .ip2(\cache_data_B[2][39] ), .op(n10511) );
  nand2_1 U13345 ( .ip1(n10575), .ip2(\cache_data_B[7][39] ), .op(n10510) );
  nand4_1 U13346 ( .ip1(n10513), .ip2(n10512), .ip3(n10511), .ip4(n10510), 
        .op(n10514) );
  not_ab_or_c_or_d U13347 ( .ip1(\cache_data_B[6][39] ), .ip2(n12337), .ip3(
        n10515), .ip4(n10514), .op(n10517) );
  nand2_1 U13348 ( .ip1(n12054), .ip2(\cache_data_B[4][39] ), .op(n10516) );
  nand3_1 U13349 ( .ip1(n10518), .ip2(n10517), .ip3(n10516), .op(n12731) );
  nand2_1 U13350 ( .ip1(n12563), .ip2(n12731), .op(n10529) );
  nand2_1 U13351 ( .ip1(n12096), .ip2(\cache_data_B[3][71] ), .op(n10527) );
  and2_1 U13352 ( .ip1(n12584), .ip2(\cache_data_B[4][71] ), .op(n10524) );
  nand2_1 U13353 ( .ip1(n11236), .ip2(\cache_data_B[5][71] ), .op(n10522) );
  nand2_1 U13354 ( .ip1(n11071), .ip2(\cache_data_B[0][71] ), .op(n10521) );
  nand2_1 U13355 ( .ip1(n10575), .ip2(\cache_data_B[7][71] ), .op(n10520) );
  nand2_1 U13356 ( .ip1(n12320), .ip2(\cache_data_B[6][71] ), .op(n10519) );
  nand4_1 U13357 ( .ip1(n10522), .ip2(n10521), .ip3(n10520), .ip4(n10519), 
        .op(n10523) );
  not_ab_or_c_or_d U13358 ( .ip1(\cache_data_B[2][71] ), .ip2(n12546), .ip3(
        n10524), .ip4(n10523), .op(n10526) );
  nand2_1 U13359 ( .ip1(n10686), .ip2(\cache_data_B[1][71] ), .op(n10525) );
  nand3_1 U13360 ( .ip1(n10527), .ip2(n10526), .ip3(n10525), .op(n12741) );
  nand2_1 U13361 ( .ip1(n12580), .ip2(n12741), .op(n10528) );
  nand4_1 U13362 ( .ip1(n10531), .ip2(n10530), .ip3(n10529), .ip4(n10528), 
        .op(n10532) );
  not_ab_or_c_or_d U13363 ( .ip1(n12550), .ip2(n12728), .ip3(n10533), .ip4(
        n10532), .op(n10544) );
  nand2_1 U13364 ( .ip1(\cache_data_B[0][103] ), .ip2(n12204), .op(n10542) );
  and2_1 U13365 ( .ip1(n12320), .ip2(\cache_data_B[6][103] ), .op(n10539) );
  nand2_1 U13366 ( .ip1(n12096), .ip2(\cache_data_B[3][103] ), .op(n10537) );
  nand2_1 U13367 ( .ip1(n10686), .ip2(\cache_data_B[1][103] ), .op(n10536) );
  nand2_1 U13368 ( .ip1(n10575), .ip2(\cache_data_B[7][103] ), .op(n10535) );
  nand2_1 U13369 ( .ip1(n11296), .ip2(\cache_data_B[5][103] ), .op(n10534) );
  nand4_1 U13370 ( .ip1(n10537), .ip2(n10536), .ip3(n10535), .ip4(n10534), 
        .op(n10538) );
  not_ab_or_c_or_d U13371 ( .ip1(n12475), .ip2(\cache_data_B[2][103] ), .ip3(
        n10539), .ip4(n10538), .op(n10541) );
  nand2_1 U13372 ( .ip1(n12054), .ip2(\cache_data_B[4][103] ), .op(n10540) );
  nand3_1 U13373 ( .ip1(n10542), .ip2(n10541), .ip3(n10540), .op(n12733) );
  nand2_1 U13374 ( .ip1(n12573), .ip2(n12733), .op(n10543) );
  nand3_1 U13375 ( .ip1(n10545), .ip2(n10544), .ip3(n10543), .op(n10546) );
  mux2_1 U13376 ( .ip1(N4183), .ip2(n10546), .s(n11472), .op(n5313) );
  nand2_1 U13377 ( .ip1(n11142), .ip2(\cache_data_A[2][104] ), .op(n10555) );
  and2_1 U13378 ( .ip1(n12147), .ip2(\cache_data_A[1][104] ), .op(n10552) );
  nand2_1 U13379 ( .ip1(n12320), .ip2(\cache_data_A[6][104] ), .op(n10550) );
  nand2_1 U13380 ( .ip1(n11071), .ip2(\cache_data_A[0][104] ), .op(n10549) );
  nand2_1 U13381 ( .ip1(n11296), .ip2(\cache_data_A[5][104] ), .op(n10548) );
  nand2_1 U13382 ( .ip1(n10575), .ip2(\cache_data_A[7][104] ), .op(n10547) );
  nand4_1 U13383 ( .ip1(n10550), .ip2(n10549), .ip3(n10548), .ip4(n10547), 
        .op(n10551) );
  not_ab_or_c_or_d U13384 ( .ip1(n11156), .ip2(\cache_data_A[4][104] ), .ip3(
        n10552), .ip4(n10551), .op(n10554) );
  nand2_1 U13385 ( .ip1(n11535), .ip2(\cache_data_A[3][104] ), .op(n10553) );
  nand3_1 U13386 ( .ip1(n10555), .ip2(n10554), .ip3(n10553), .op(n12748) );
  nand2_1 U13387 ( .ip1(n12509), .ip2(n12748), .op(n10629) );
  nand2_1 U13388 ( .ip1(n11071), .ip2(\cache_data_A[0][8] ), .op(n10564) );
  and2_1 U13389 ( .ip1(n10686), .ip2(\cache_data_A[1][8] ), .op(n10561) );
  nand2_1 U13390 ( .ip1(n12054), .ip2(\cache_data_A[4][8] ), .op(n10559) );
  nand2_1 U13391 ( .ip1(n11142), .ip2(\cache_data_A[2][8] ), .op(n10558) );
  nand2_1 U13392 ( .ip1(n11236), .ip2(\cache_data_A[5][8] ), .op(n10557) );
  nand2_1 U13393 ( .ip1(n11780), .ip2(\cache_data_A[6][8] ), .op(n10556) );
  nand4_1 U13394 ( .ip1(n10559), .ip2(n10558), .ip3(n10557), .ip4(n10556), 
        .op(n10560) );
  not_ab_or_c_or_d U13395 ( .ip1(\cache_data_A[7][8] ), .ip2(n12278), .ip3(
        n10561), .ip4(n10560), .op(n10563) );
  nand2_1 U13396 ( .ip1(n12096), .ip2(\cache_data_A[3][8] ), .op(n10562) );
  nand3_1 U13397 ( .ip1(n10564), .ip2(n10563), .ip3(n10562), .op(n12749) );
  nand2_1 U13398 ( .ip1(n12054), .ip2(\cache_data_A[4][72] ), .op(n10568) );
  nand2_1 U13399 ( .ip1(n11071), .ip2(\cache_data_A[0][72] ), .op(n10567) );
  nand2_1 U13400 ( .ip1(n11142), .ip2(\cache_data_A[2][72] ), .op(n10566) );
  nand2_1 U13401 ( .ip1(n10575), .ip2(\cache_data_A[7][72] ), .op(n10565) );
  nand4_1 U13402 ( .ip1(n10568), .ip2(n10567), .ip3(n10566), .ip4(n10565), 
        .op(n10574) );
  nand2_1 U13403 ( .ip1(n12337), .ip2(\cache_data_A[6][72] ), .op(n10572) );
  nand2_1 U13404 ( .ip1(n11724), .ip2(\cache_data_A[1][72] ), .op(n10571) );
  nand2_1 U13405 ( .ip1(n11236), .ip2(\cache_data_A[5][72] ), .op(n10570) );
  nand2_1 U13406 ( .ip1(n12559), .ip2(\cache_data_A[3][72] ), .op(n10569) );
  nand4_1 U13407 ( .ip1(n10572), .ip2(n10571), .ip3(n10570), .ip4(n10569), 
        .op(n10573) );
  nor2_1 U13408 ( .ip1(n10574), .ip2(n10573), .op(n12747) );
  nor2_1 U13409 ( .ip1(n12747), .ip2(n12529), .op(n10617) );
  nand2_1 U13410 ( .ip1(\cache_data_B[3][104] ), .ip2(n12410), .op(n10584) );
  and2_1 U13411 ( .ip1(n12486), .ip2(\cache_data_B[2][104] ), .op(n10581) );
  nand2_1 U13412 ( .ip1(n12054), .ip2(\cache_data_B[4][104] ), .op(n10579) );
  nand2_1 U13413 ( .ip1(n12337), .ip2(\cache_data_B[6][104] ), .op(n10578) );
  nand2_1 U13414 ( .ip1(n11304), .ip2(\cache_data_B[5][104] ), .op(n10577) );
  nand2_1 U13415 ( .ip1(n10575), .ip2(\cache_data_B[7][104] ), .op(n10576) );
  nand4_1 U13416 ( .ip1(n10579), .ip2(n10578), .ip3(n10577), .ip4(n10576), 
        .op(n10580) );
  not_ab_or_c_or_d U13417 ( .ip1(\cache_data_B[0][104] ), .ip2(n12297), .ip3(
        n10581), .ip4(n10580), .op(n10583) );
  nand2_1 U13418 ( .ip1(n11724), .ip2(\cache_data_B[1][104] ), .op(n10582) );
  nand3_1 U13419 ( .ip1(n10584), .ip2(n10583), .ip3(n10582), .op(n12758) );
  nand2_1 U13420 ( .ip1(n12573), .ip2(n12758), .op(n10615) );
  nand2_1 U13421 ( .ip1(n12337), .ip2(\cache_data_B[6][72] ), .op(n10593) );
  and2_1 U13422 ( .ip1(n12582), .ip2(\cache_data_B[5][72] ), .op(n10590) );
  nand2_1 U13423 ( .ip1(n11071), .ip2(\cache_data_B[0][72] ), .op(n10588) );
  nand2_1 U13424 ( .ip1(n11535), .ip2(\cache_data_B[3][72] ), .op(n10587) );
  nand2_1 U13425 ( .ip1(n11142), .ip2(\cache_data_B[2][72] ), .op(n10586) );
  nand2_1 U13426 ( .ip1(n10686), .ip2(\cache_data_B[1][72] ), .op(n10585) );
  nand4_1 U13427 ( .ip1(n10588), .ip2(n10587), .ip3(n10586), .ip4(n10585), 
        .op(n10589) );
  not_ab_or_c_or_d U13428 ( .ip1(\cache_data_B[7][72] ), .ip2(n12278), .ip3(
        n10590), .ip4(n10589), .op(n10592) );
  nand2_1 U13429 ( .ip1(n12054), .ip2(\cache_data_B[4][72] ), .op(n10591) );
  nand3_1 U13430 ( .ip1(n10593), .ip2(n10592), .ip3(n10591), .op(n12751) );
  nand2_1 U13431 ( .ip1(n12580), .ip2(n12751), .op(n10614) );
  nand2_1 U13432 ( .ip1(n10702), .ip2(\cache_data_B[7][40] ), .op(n10602) );
  and2_1 U13433 ( .ip1(n12458), .ip2(\cache_data_B[6][40] ), .op(n10599) );
  nand2_1 U13434 ( .ip1(n11280), .ip2(\cache_data_B[5][40] ), .op(n10597) );
  nand2_1 U13435 ( .ip1(n11071), .ip2(\cache_data_B[0][40] ), .op(n10596) );
  nand2_1 U13436 ( .ip1(n12054), .ip2(\cache_data_B[4][40] ), .op(n10595) );
  nand2_1 U13437 ( .ip1(n11724), .ip2(\cache_data_B[1][40] ), .op(n10594) );
  nand4_1 U13438 ( .ip1(n10597), .ip2(n10596), .ip3(n10595), .ip4(n10594), 
        .op(n10598) );
  not_ab_or_c_or_d U13439 ( .ip1(n12546), .ip2(\cache_data_B[2][40] ), .ip3(
        n10599), .ip4(n10598), .op(n10601) );
  nand2_1 U13440 ( .ip1(n12096), .ip2(\cache_data_B[3][40] ), .op(n10600) );
  nand3_1 U13441 ( .ip1(n10602), .ip2(n10601), .ip3(n10600), .op(n12759) );
  nand2_1 U13442 ( .ip1(n12563), .ip2(n12759), .op(n10613) );
  nand2_1 U13443 ( .ip1(\cache_data_A[6][40] ), .ip2(n12458), .op(n10611) );
  and2_1 U13444 ( .ip1(n12147), .ip2(\cache_data_A[1][40] ), .op(n10608) );
  nand2_1 U13445 ( .ip1(n12096), .ip2(\cache_data_A[3][40] ), .op(n10606) );
  nand2_1 U13446 ( .ip1(n10702), .ip2(\cache_data_A[7][40] ), .op(n10605) );
  nand2_1 U13447 ( .ip1(n11236), .ip2(\cache_data_A[5][40] ), .op(n10604) );
  nand2_1 U13448 ( .ip1(n11071), .ip2(\cache_data_A[0][40] ), .op(n10603) );
  nand4_1 U13449 ( .ip1(n10606), .ip2(n10605), .ip3(n10604), .ip4(n10603), 
        .op(n10607) );
  not_ab_or_c_or_d U13450 ( .ip1(n12546), .ip2(\cache_data_A[2][40] ), .ip3(
        n10608), .ip4(n10607), .op(n10610) );
  nand2_1 U13451 ( .ip1(n12054), .ip2(\cache_data_A[4][40] ), .op(n10609) );
  nand3_1 U13452 ( .ip1(n10611), .ip2(n10610), .ip3(n10609), .op(n12750) );
  nand2_1 U13453 ( .ip1(n12595), .ip2(n12750), .op(n10612) );
  nand4_1 U13454 ( .ip1(n10615), .ip2(n10614), .ip3(n10613), .ip4(n10612), 
        .op(n10616) );
  not_ab_or_c_or_d U13455 ( .ip1(n12550), .ip2(n12749), .ip3(n10617), .ip4(
        n10616), .op(n10628) );
  nand2_1 U13456 ( .ip1(n11071), .ip2(\cache_data_B[0][8] ), .op(n10626) );
  and2_1 U13457 ( .ip1(n12410), .ip2(\cache_data_B[3][8] ), .op(n10623) );
  nand2_1 U13458 ( .ip1(n11280), .ip2(\cache_data_B[5][8] ), .op(n10621) );
  nand2_1 U13459 ( .ip1(n11142), .ip2(\cache_data_B[2][8] ), .op(n10620) );
  nand2_1 U13460 ( .ip1(n12054), .ip2(\cache_data_B[4][8] ), .op(n10619) );
  nand2_1 U13461 ( .ip1(n11724), .ip2(\cache_data_B[1][8] ), .op(n10618) );
  nand4_1 U13462 ( .ip1(n10621), .ip2(n10620), .ip3(n10619), .ip4(n10618), 
        .op(n10622) );
  not_ab_or_c_or_d U13463 ( .ip1(\cache_data_B[7][8] ), .ip2(n12278), .ip3(
        n10623), .ip4(n10622), .op(n10625) );
  nand2_1 U13464 ( .ip1(n12337), .ip2(\cache_data_B[6][8] ), .op(n10624) );
  nand3_1 U13465 ( .ip1(n10626), .ip2(n10625), .ip3(n10624), .op(n12746) );
  nand2_1 U13466 ( .ip1(n12539), .ip2(n12746), .op(n10627) );
  nand3_1 U13467 ( .ip1(n10629), .ip2(n10628), .ip3(n10627), .op(n10630) );
  mux2_1 U13468 ( .ip1(N4180), .ip2(n10630), .s(n11472), .op(n5312) );
  nand2_1 U13469 ( .ip1(n11142), .ip2(\cache_data_A[2][105] ), .op(n10639) );
  and2_1 U13470 ( .ip1(n12371), .ip2(\cache_data_A[6][105] ), .op(n10636) );
  nand2_1 U13471 ( .ip1(n12559), .ip2(\cache_data_A[3][105] ), .op(n10634) );
  nand2_1 U13472 ( .ip1(n11071), .ip2(\cache_data_A[0][105] ), .op(n10633) );
  nand2_1 U13473 ( .ip1(n11236), .ip2(\cache_data_A[5][105] ), .op(n10632) );
  nand2_1 U13474 ( .ip1(n10686), .ip2(\cache_data_A[1][105] ), .op(n10631) );
  nand4_1 U13475 ( .ip1(n10634), .ip2(n10633), .ip3(n10632), .ip4(n10631), 
        .op(n10635) );
  not_ab_or_c_or_d U13476 ( .ip1(\cache_data_A[7][105] ), .ip2(n11057), .ip3(
        n10636), .ip4(n10635), .op(n10638) );
  nand2_1 U13477 ( .ip1(n11324), .ip2(\cache_data_A[4][105] ), .op(n10637) );
  nand3_1 U13478 ( .ip1(n10639), .ip2(n10638), .ip3(n10637), .op(n12777) );
  nand2_1 U13479 ( .ip1(n12509), .ip2(n12777), .op(n10714) );
  nand2_1 U13480 ( .ip1(n11071), .ip2(\cache_data_B[0][9] ), .op(n10648) );
  and2_1 U13481 ( .ip1(n12194), .ip2(\cache_data_B[4][9] ), .op(n10645) );
  nand2_1 U13482 ( .ip1(n10702), .ip2(\cache_data_B[7][9] ), .op(n10643) );
  nand2_1 U13483 ( .ip1(n11535), .ip2(\cache_data_B[3][9] ), .op(n10642) );
  nand2_1 U13484 ( .ip1(n12337), .ip2(\cache_data_B[6][9] ), .op(n10641) );
  nand2_1 U13485 ( .ip1(n11280), .ip2(\cache_data_B[5][9] ), .op(n10640) );
  nand4_1 U13486 ( .ip1(n10643), .ip2(n10642), .ip3(n10641), .ip4(n10640), 
        .op(n10644) );
  not_ab_or_c_or_d U13487 ( .ip1(n12546), .ip2(\cache_data_B[2][9] ), .ip3(
        n10645), .ip4(n10644), .op(n10647) );
  nand2_1 U13488 ( .ip1(n11724), .ip2(\cache_data_B[1][9] ), .op(n10646) );
  nand3_1 U13489 ( .ip1(n10648), .ip2(n10647), .ip3(n10646), .op(n12768) );
  nand2_1 U13490 ( .ip1(n11304), .ip2(\cache_data_A[5][73] ), .op(n10652) );
  nand2_1 U13491 ( .ip1(n12337), .ip2(\cache_data_A[6][73] ), .op(n10651) );
  nand2_1 U13492 ( .ip1(n11724), .ip2(\cache_data_A[1][73] ), .op(n10650) );
  nand2_1 U13493 ( .ip1(n12357), .ip2(\cache_data_A[0][73] ), .op(n10649) );
  nand4_1 U13494 ( .ip1(n10652), .ip2(n10651), .ip3(n10650), .ip4(n10649), 
        .op(n10658) );
  nand2_1 U13495 ( .ip1(n12096), .ip2(\cache_data_A[3][73] ), .op(n10656) );
  nand2_1 U13496 ( .ip1(n11156), .ip2(\cache_data_A[4][73] ), .op(n10655) );
  nand2_1 U13497 ( .ip1(n10702), .ip2(\cache_data_A[7][73] ), .op(n10654) );
  nand2_1 U13498 ( .ip1(n11142), .ip2(\cache_data_A[2][73] ), .op(n10653) );
  nand4_1 U13499 ( .ip1(n10656), .ip2(n10655), .ip3(n10654), .ip4(n10653), 
        .op(n10657) );
  nor2_1 U13500 ( .ip1(n10658), .ip2(n10657), .op(n12765) );
  nor2_1 U13501 ( .ip1(n12765), .ip2(n12529), .op(n10701) );
  nand2_1 U13502 ( .ip1(\cache_data_A[3][41] ), .ip2(n12410), .op(n10667) );
  and2_1 U13503 ( .ip1(n12486), .ip2(\cache_data_A[2][41] ), .op(n10664) );
  nand2_1 U13504 ( .ip1(n12337), .ip2(\cache_data_A[6][41] ), .op(n10662) );
  nand2_1 U13505 ( .ip1(n10702), .ip2(\cache_data_A[7][41] ), .op(n10661) );
  nand2_1 U13506 ( .ip1(n11236), .ip2(\cache_data_A[5][41] ), .op(n10660) );
  nand2_1 U13507 ( .ip1(n11156), .ip2(\cache_data_A[4][41] ), .op(n10659) );
  nand4_1 U13508 ( .ip1(n10662), .ip2(n10661), .ip3(n10660), .ip4(n10659), 
        .op(n10663) );
  not_ab_or_c_or_d U13509 ( .ip1(\cache_data_A[0][41] ), .ip2(n12297), .ip3(
        n10664), .ip4(n10663), .op(n10666) );
  nand2_1 U13510 ( .ip1(n10686), .ip2(\cache_data_A[1][41] ), .op(n10665) );
  nand3_1 U13511 ( .ip1(n10667), .ip2(n10666), .ip3(n10665), .op(n12767) );
  nand2_1 U13512 ( .ip1(n12595), .ip2(n12767), .op(n10699) );
  nand2_1 U13513 ( .ip1(n12337), .ip2(\cache_data_B[6][105] ), .op(n10676) );
  and2_1 U13514 ( .ip1(n12147), .ip2(\cache_data_B[1][105] ), .op(n10673) );
  nand2_1 U13515 ( .ip1(n12357), .ip2(\cache_data_B[0][105] ), .op(n10671) );
  nand2_1 U13516 ( .ip1(n12054), .ip2(\cache_data_B[4][105] ), .op(n10670) );
  nand2_1 U13517 ( .ip1(n11280), .ip2(\cache_data_B[5][105] ), .op(n10669) );
  nand2_1 U13518 ( .ip1(n11142), .ip2(\cache_data_B[2][105] ), .op(n10668) );
  nand4_1 U13519 ( .ip1(n10671), .ip2(n10670), .ip3(n10669), .ip4(n10668), 
        .op(n10672) );
  not_ab_or_c_or_d U13520 ( .ip1(n12278), .ip2(\cache_data_B[7][105] ), .ip3(
        n10673), .ip4(n10672), .op(n10675) );
  nand2_1 U13521 ( .ip1(n11535), .ip2(\cache_data_B[3][105] ), .op(n10674) );
  nand3_1 U13522 ( .ip1(n10676), .ip2(n10675), .ip3(n10674), .op(n12776) );
  nand2_1 U13523 ( .ip1(n12573), .ip2(n12776), .op(n10698) );
  nand2_1 U13524 ( .ip1(\cache_data_B[0][73] ), .ip2(n12204), .op(n10685) );
  and2_1 U13525 ( .ip1(n12396), .ip2(\cache_data_B[4][73] ), .op(n10682) );
  nand2_1 U13526 ( .ip1(n11142), .ip2(\cache_data_B[2][73] ), .op(n10680) );
  nand2_1 U13527 ( .ip1(n10686), .ip2(\cache_data_B[1][73] ), .op(n10679) );
  nand2_1 U13528 ( .ip1(n11236), .ip2(\cache_data_B[5][73] ), .op(n10678) );
  nand2_1 U13529 ( .ip1(n11535), .ip2(\cache_data_B[3][73] ), .op(n10677) );
  nand4_1 U13530 ( .ip1(n10680), .ip2(n10679), .ip3(n10678), .ip4(n10677), 
        .op(n10681) );
  not_ab_or_c_or_d U13531 ( .ip1(\cache_data_B[6][73] ), .ip2(n12337), .ip3(
        n10682), .ip4(n10681), .op(n10684) );
  nand2_1 U13532 ( .ip1(n10702), .ip2(\cache_data_B[7][73] ), .op(n10683) );
  nand3_1 U13533 ( .ip1(n10685), .ip2(n10684), .ip3(n10683), .op(n12769) );
  nand2_1 U13534 ( .ip1(n12580), .ip2(n12769), .op(n10697) );
  nand2_1 U13535 ( .ip1(\cache_data_B[2][41] ), .ip2(n12486), .op(n10695) );
  and2_1 U13536 ( .ip1(n12256), .ip2(\cache_data_B[5][41] ), .op(n10692) );
  nand2_1 U13537 ( .ip1(n10686), .ip2(\cache_data_B[1][41] ), .op(n10690) );
  nand2_1 U13538 ( .ip1(n11535), .ip2(\cache_data_B[3][41] ), .op(n10689) );
  nand2_1 U13539 ( .ip1(n12337), .ip2(\cache_data_B[6][41] ), .op(n10688) );
  nand2_1 U13540 ( .ip1(n10702), .ip2(\cache_data_B[7][41] ), .op(n10687) );
  nand4_1 U13541 ( .ip1(n10690), .ip2(n10689), .ip3(n10688), .ip4(n10687), 
        .op(n10691) );
  not_ab_or_c_or_d U13542 ( .ip1(n12297), .ip2(\cache_data_B[0][41] ), .ip3(
        n10692), .ip4(n10691), .op(n10694) );
  nand2_1 U13543 ( .ip1(n11156), .ip2(\cache_data_B[4][41] ), .op(n10693) );
  nand3_1 U13544 ( .ip1(n10695), .ip2(n10694), .ip3(n10693), .op(n12766) );
  nand2_1 U13545 ( .ip1(n12563), .ip2(n12766), .op(n10696) );
  nand4_1 U13546 ( .ip1(n10699), .ip2(n10698), .ip3(n10697), .ip4(n10696), 
        .op(n10700) );
  not_ab_or_c_or_d U13547 ( .ip1(n12539), .ip2(n12768), .ip3(n10701), .ip4(
        n10700), .op(n10713) );
  nand2_1 U13548 ( .ip1(n10702), .ip2(\cache_data_A[7][9] ), .op(n10711) );
  and2_1 U13549 ( .ip1(n11296), .ip2(\cache_data_A[5][9] ), .op(n10708) );
  nand2_1 U13550 ( .ip1(n12559), .ip2(\cache_data_A[3][9] ), .op(n10706) );
  nand2_1 U13551 ( .ip1(n11071), .ip2(\cache_data_A[0][9] ), .op(n10705) );
  nand2_1 U13552 ( .ip1(n11324), .ip2(\cache_data_A[4][9] ), .op(n10704) );
  nand2_1 U13553 ( .ip1(n12337), .ip2(\cache_data_A[6][9] ), .op(n10703) );
  nand4_1 U13554 ( .ip1(n10706), .ip2(n10705), .ip3(n10704), .ip4(n10703), 
        .op(n10707) );
  not_ab_or_c_or_d U13555 ( .ip1(\cache_data_A[2][9] ), .ip2(n12546), .ip3(
        n10708), .ip4(n10707), .op(n10710) );
  nand2_1 U13556 ( .ip1(n11724), .ip2(\cache_data_A[1][9] ), .op(n10709) );
  nand3_1 U13557 ( .ip1(n10711), .ip2(n10710), .ip3(n10709), .op(n12764) );
  nand2_1 U13558 ( .ip1(n12550), .ip2(n12764), .op(n10712) );
  nand3_1 U13559 ( .ip1(n10714), .ip2(n10713), .ip3(n10712), .op(n10715) );
  mux2_1 U13560 ( .ip1(N4177), .ip2(n10715), .s(n11472), .op(n5311) );
  nand2_1 U13561 ( .ip1(\cache_data_B[2][106] ), .ip2(n12486), .op(n10724) );
  and2_1 U13562 ( .ip1(n12194), .ip2(\cache_data_B[4][106] ), .op(n10721) );
  nand2_1 U13563 ( .ip1(n11535), .ip2(\cache_data_B[3][106] ), .op(n10719) );
  nand2_1 U13564 ( .ip1(n11057), .ip2(\cache_data_B[7][106] ), .op(n10718) );
  nand2_1 U13565 ( .ip1(n12337), .ip2(\cache_data_B[6][106] ), .op(n10717) );
  buf_1 U13566 ( .ip(n11724), .op(n11311) );
  nand2_1 U13567 ( .ip1(n11311), .ip2(\cache_data_B[1][106] ), .op(n10716) );
  nand4_1 U13568 ( .ip1(n10719), .ip2(n10718), .ip3(n10717), .ip4(n10716), 
        .op(n10720) );
  not_ab_or_c_or_d U13569 ( .ip1(\cache_data_B[0][106] ), .ip2(n12297), .ip3(
        n10721), .ip4(n10720), .op(n10723) );
  nand2_1 U13570 ( .ip1(n11304), .ip2(\cache_data_B[5][106] ), .op(n10722) );
  nand3_1 U13571 ( .ip1(n10724), .ip2(n10723), .ip3(n10722), .op(n12786) );
  nand2_1 U13572 ( .ip1(n12573), .ip2(n12786), .op(n10797) );
  nand2_1 U13573 ( .ip1(\cache_data_B[7][42] ), .ip2(n12552), .op(n10733) );
  and2_1 U13574 ( .ip1(n10686), .ip2(\cache_data_B[1][42] ), .op(n10730) );
  nand2_1 U13575 ( .ip1(n11535), .ip2(\cache_data_B[3][42] ), .op(n10728) );
  nand2_1 U13576 ( .ip1(n12337), .ip2(\cache_data_B[6][42] ), .op(n10727) );
  nand2_1 U13577 ( .ip1(n12357), .ip2(\cache_data_B[0][42] ), .op(n10726) );
  nand2_1 U13578 ( .ip1(n12584), .ip2(\cache_data_B[4][42] ), .op(n10725) );
  nand4_1 U13579 ( .ip1(n10728), .ip2(n10727), .ip3(n10726), .ip4(n10725), 
        .op(n10729) );
  not_ab_or_c_or_d U13580 ( .ip1(n12546), .ip2(\cache_data_B[2][42] ), .ip3(
        n10730), .ip4(n10729), .op(n10732) );
  nand2_1 U13581 ( .ip1(n11304), .ip2(\cache_data_B[5][42] ), .op(n10731) );
  nand3_1 U13582 ( .ip1(n10733), .ip2(n10732), .ip3(n10731), .op(n12787) );
  nand2_1 U13583 ( .ip1(n11311), .ip2(\cache_data_A[1][74] ), .op(n10737) );
  nand2_1 U13584 ( .ip1(n11304), .ip2(\cache_data_A[5][74] ), .op(n10736) );
  nand2_1 U13585 ( .ip1(n11142), .ip2(\cache_data_A[2][74] ), .op(n10735) );
  nand2_1 U13586 ( .ip1(n11057), .ip2(\cache_data_A[7][74] ), .op(n10734) );
  nand4_1 U13587 ( .ip1(n10737), .ip2(n10736), .ip3(n10735), .ip4(n10734), 
        .op(n10743) );
  nand2_1 U13588 ( .ip1(n12559), .ip2(\cache_data_A[3][74] ), .op(n10741) );
  nand2_1 U13589 ( .ip1(n12337), .ip2(\cache_data_A[6][74] ), .op(n10740) );
  nand2_1 U13590 ( .ip1(n12357), .ip2(\cache_data_A[0][74] ), .op(n10739) );
  nand2_1 U13591 ( .ip1(n11324), .ip2(\cache_data_A[4][74] ), .op(n10738) );
  nand4_1 U13592 ( .ip1(n10741), .ip2(n10740), .ip3(n10739), .ip4(n10738), 
        .op(n10742) );
  nor2_1 U13593 ( .ip1(n10743), .ip2(n10742), .op(n12783) );
  nor2_1 U13594 ( .ip1(n12783), .ip2(n12529), .op(n10785) );
  nand2_1 U13595 ( .ip1(n12357), .ip2(\cache_data_A[0][42] ), .op(n10752) );
  and2_1 U13596 ( .ip1(n12194), .ip2(\cache_data_A[4][42] ), .op(n10749) );
  nand2_1 U13597 ( .ip1(n11304), .ip2(\cache_data_A[5][42] ), .op(n10747) );
  nand2_1 U13598 ( .ip1(n11311), .ip2(\cache_data_A[1][42] ), .op(n10746) );
  nand2_1 U13599 ( .ip1(n12320), .ip2(\cache_data_A[6][42] ), .op(n10745) );
  nand2_1 U13600 ( .ip1(n11142), .ip2(\cache_data_A[2][42] ), .op(n10744) );
  nand4_1 U13601 ( .ip1(n10747), .ip2(n10746), .ip3(n10745), .ip4(n10744), 
        .op(n10748) );
  not_ab_or_c_or_d U13602 ( .ip1(\cache_data_A[7][42] ), .ip2(n12278), .ip3(
        n10749), .ip4(n10748), .op(n10751) );
  nand2_1 U13603 ( .ip1(n12559), .ip2(\cache_data_A[3][42] ), .op(n10750) );
  nand3_1 U13604 ( .ip1(n10752), .ip2(n10751), .ip3(n10750), .op(n12795) );
  nand2_1 U13605 ( .ip1(n12595), .ip2(n12795), .op(n10783) );
  nand2_1 U13606 ( .ip1(n11142), .ip2(\cache_data_B[2][74] ), .op(n10761) );
  and2_1 U13607 ( .ip1(n10686), .ip2(\cache_data_B[1][74] ), .op(n10758) );
  nand2_1 U13608 ( .ip1(n12320), .ip2(\cache_data_B[6][74] ), .op(n10756) );
  nand2_1 U13609 ( .ip1(n11071), .ip2(\cache_data_B[0][74] ), .op(n10755) );
  nand2_1 U13610 ( .ip1(n11296), .ip2(\cache_data_B[5][74] ), .op(n10754) );
  nand2_1 U13611 ( .ip1(n12054), .ip2(\cache_data_B[4][74] ), .op(n10753) );
  nand4_1 U13612 ( .ip1(n10756), .ip2(n10755), .ip3(n10754), .ip4(n10753), 
        .op(n10757) );
  not_ab_or_c_or_d U13613 ( .ip1(\cache_data_B[3][74] ), .ip2(n11535), .ip3(
        n10758), .ip4(n10757), .op(n10760) );
  nand2_1 U13614 ( .ip1(n11057), .ip2(\cache_data_B[7][74] ), .op(n10759) );
  nand3_1 U13615 ( .ip1(n10761), .ip2(n10760), .ip3(n10759), .op(n12794) );
  nand2_1 U13616 ( .ip1(n12580), .ip2(n12794), .op(n10782) );
  nand2_1 U13617 ( .ip1(n11142), .ip2(\cache_data_A[2][10] ), .op(n10770) );
  and2_1 U13618 ( .ip1(n12147), .ip2(\cache_data_A[1][10] ), .op(n10767) );
  nand2_1 U13619 ( .ip1(n12320), .ip2(\cache_data_A[6][10] ), .op(n10765) );
  nand2_1 U13620 ( .ip1(n12357), .ip2(\cache_data_A[0][10] ), .op(n10764) );
  nand2_1 U13621 ( .ip1(n11057), .ip2(\cache_data_A[7][10] ), .op(n10763) );
  nand2_1 U13622 ( .ip1(n11304), .ip2(\cache_data_A[5][10] ), .op(n10762) );
  nand4_1 U13623 ( .ip1(n10765), .ip2(n10764), .ip3(n10763), .ip4(n10762), 
        .op(n10766) );
  not_ab_or_c_or_d U13624 ( .ip1(\cache_data_A[3][10] ), .ip2(n12559), .ip3(
        n10767), .ip4(n10766), .op(n10769) );
  nand2_1 U13625 ( .ip1(n12476), .ip2(\cache_data_A[4][10] ), .op(n10768) );
  nand3_1 U13626 ( .ip1(n10770), .ip2(n10769), .ip3(n10768), .op(n12785) );
  nand2_1 U13627 ( .ip1(n12550), .ip2(n12785), .op(n10781) );
  nand2_1 U13628 ( .ip1(n11142), .ip2(\cache_data_A[2][106] ), .op(n10779) );
  and2_1 U13629 ( .ip1(n12582), .ip2(\cache_data_A[5][106] ), .op(n10776) );
  nand2_1 U13630 ( .ip1(n11311), .ip2(\cache_data_A[1][106] ), .op(n10774) );
  nand2_1 U13631 ( .ip1(n11535), .ip2(\cache_data_A[3][106] ), .op(n10773) );
  nand2_1 U13632 ( .ip1(n11057), .ip2(\cache_data_A[7][106] ), .op(n10772) );
  nand2_1 U13633 ( .ip1(n12357), .ip2(\cache_data_A[0][106] ), .op(n10771) );
  nand4_1 U13634 ( .ip1(n10774), .ip2(n10773), .ip3(n10772), .ip4(n10771), 
        .op(n10775) );
  not_ab_or_c_or_d U13635 ( .ip1(\cache_data_A[6][106] ), .ip2(n12337), .ip3(
        n10776), .ip4(n10775), .op(n10778) );
  nand2_1 U13636 ( .ip1(n12054), .ip2(\cache_data_A[4][106] ), .op(n10777) );
  nand3_1 U13637 ( .ip1(n10779), .ip2(n10778), .ip3(n10777), .op(n12784) );
  nand2_1 U13638 ( .ip1(n12509), .ip2(n12784), .op(n10780) );
  nand4_1 U13639 ( .ip1(n10783), .ip2(n10782), .ip3(n10781), .ip4(n10780), 
        .op(n10784) );
  not_ab_or_c_or_d U13640 ( .ip1(n12563), .ip2(n12787), .ip3(n10785), .ip4(
        n10784), .op(n10796) );
  nand2_1 U13641 ( .ip1(n12559), .ip2(\cache_data_B[3][10] ), .op(n10794) );
  and2_1 U13642 ( .ip1(n12476), .ip2(\cache_data_B[4][10] ), .op(n10791) );
  nand2_1 U13643 ( .ip1(n11236), .ip2(\cache_data_B[5][10] ), .op(n10789) );
  nand2_1 U13644 ( .ip1(n11142), .ip2(\cache_data_B[2][10] ), .op(n10788) );
  nand2_1 U13645 ( .ip1(n12357), .ip2(\cache_data_B[0][10] ), .op(n10787) );
  nand2_1 U13646 ( .ip1(n11057), .ip2(\cache_data_B[7][10] ), .op(n10786) );
  nand4_1 U13647 ( .ip1(n10789), .ip2(n10788), .ip3(n10787), .ip4(n10786), 
        .op(n10790) );
  not_ab_or_c_or_d U13648 ( .ip1(n12551), .ip2(\cache_data_B[6][10] ), .ip3(
        n10791), .ip4(n10790), .op(n10793) );
  nand2_1 U13649 ( .ip1(n11311), .ip2(\cache_data_B[1][10] ), .op(n10792) );
  nand3_1 U13650 ( .ip1(n10794), .ip2(n10793), .ip3(n10792), .op(n12782) );
  nand2_1 U13651 ( .ip1(n12539), .ip2(n12782), .op(n10795) );
  nand3_1 U13652 ( .ip1(n10797), .ip2(n10796), .ip3(n10795), .op(n10798) );
  mux2_1 U13653 ( .ip1(N4174), .ip2(n10798), .s(n11472), .op(n5310) );
  nand2_1 U13654 ( .ip1(n11535), .ip2(\cache_data_A[3][107] ), .op(n10807) );
  and2_1 U13655 ( .ip1(n12147), .ip2(\cache_data_A[1][107] ), .op(n10804) );
  nand2_1 U13656 ( .ip1(n12584), .ip2(\cache_data_A[4][107] ), .op(n10802) );
  nand2_1 U13657 ( .ip1(n11142), .ip2(\cache_data_A[2][107] ), .op(n10801) );
  nand2_1 U13658 ( .ip1(n12357), .ip2(\cache_data_A[0][107] ), .op(n10800) );
  nand2_1 U13659 ( .ip1(n12371), .ip2(\cache_data_A[6][107] ), .op(n10799) );
  nand4_1 U13660 ( .ip1(n10802), .ip2(n10801), .ip3(n10800), .ip4(n10799), 
        .op(n10803) );
  not_ab_or_c_or_d U13661 ( .ip1(n12278), .ip2(\cache_data_A[7][107] ), .ip3(
        n10804), .ip4(n10803), .op(n10806) );
  nand2_1 U13662 ( .ip1(n11304), .ip2(\cache_data_A[5][107] ), .op(n10805) );
  nand3_1 U13663 ( .ip1(n10807), .ip2(n10806), .ip3(n10805), .op(n12805) );
  nand2_1 U13664 ( .ip1(n12509), .ip2(n12805), .op(n10880) );
  nand2_1 U13665 ( .ip1(n11142), .ip2(\cache_data_A[2][11] ), .op(n10816) );
  and2_1 U13666 ( .ip1(n12476), .ip2(\cache_data_A[4][11] ), .op(n10813) );
  nand2_1 U13667 ( .ip1(n11311), .ip2(\cache_data_A[1][11] ), .op(n10811) );
  nand2_1 U13668 ( .ip1(n11280), .ip2(\cache_data_A[5][11] ), .op(n10810) );
  nand2_1 U13669 ( .ip1(n11057), .ip2(\cache_data_A[7][11] ), .op(n10809) );
  nand2_1 U13670 ( .ip1(n12357), .ip2(\cache_data_A[0][11] ), .op(n10808) );
  nand4_1 U13671 ( .ip1(n10811), .ip2(n10810), .ip3(n10809), .ip4(n10808), 
        .op(n10812) );
  not_ab_or_c_or_d U13672 ( .ip1(\cache_data_A[6][11] ), .ip2(n12337), .ip3(
        n10813), .ip4(n10812), .op(n10815) );
  nand2_1 U13673 ( .ip1(n12096), .ip2(\cache_data_A[3][11] ), .op(n10814) );
  nand3_1 U13674 ( .ip1(n10816), .ip2(n10815), .ip3(n10814), .op(n12803) );
  nand2_1 U13675 ( .ip1(n12357), .ip2(\cache_data_A[0][75] ), .op(n10820) );
  nand2_1 U13676 ( .ip1(n12468), .ip2(\cache_data_A[7][75] ), .op(n10819) );
  nand2_1 U13677 ( .ip1(n12320), .ip2(\cache_data_A[6][75] ), .op(n10818) );
  nand2_1 U13678 ( .ip1(n12559), .ip2(\cache_data_A[3][75] ), .op(n10817) );
  nand4_1 U13679 ( .ip1(n10820), .ip2(n10819), .ip3(n10818), .ip4(n10817), 
        .op(n10826) );
  nand2_1 U13680 ( .ip1(n11142), .ip2(\cache_data_A[2][75] ), .op(n10824) );
  nand2_1 U13681 ( .ip1(n11311), .ip2(\cache_data_A[1][75] ), .op(n10823) );
  nand2_1 U13682 ( .ip1(n11236), .ip2(\cache_data_A[5][75] ), .op(n10822) );
  nand2_1 U13683 ( .ip1(n11324), .ip2(\cache_data_A[4][75] ), .op(n10821) );
  nand4_1 U13684 ( .ip1(n10824), .ip2(n10823), .ip3(n10822), .ip4(n10821), 
        .op(n10825) );
  nor2_1 U13685 ( .ip1(n10826), .ip2(n10825), .op(n12801) );
  nor2_1 U13686 ( .ip1(n12801), .ip2(n12529), .op(n10868) );
  nand2_1 U13687 ( .ip1(n12357), .ip2(\cache_data_B[0][75] ), .op(n10835) );
  and2_1 U13688 ( .ip1(n8060), .ip2(\cache_data_B[3][75] ), .op(n10832) );
  nand2_1 U13689 ( .ip1(n12278), .ip2(\cache_data_B[7][75] ), .op(n10830) );
  nand2_1 U13690 ( .ip1(n12320), .ip2(\cache_data_B[6][75] ), .op(n10829) );
  nand2_1 U13691 ( .ip1(n11311), .ip2(\cache_data_B[1][75] ), .op(n10828) );
  nand2_1 U13692 ( .ip1(n11304), .ip2(\cache_data_B[5][75] ), .op(n10827) );
  nand4_1 U13693 ( .ip1(n10830), .ip2(n10829), .ip3(n10828), .ip4(n10827), 
        .op(n10831) );
  not_ab_or_c_or_d U13694 ( .ip1(\cache_data_B[2][75] ), .ip2(n12546), .ip3(
        n10832), .ip4(n10831), .op(n10834) );
  nand2_1 U13695 ( .ip1(n11324), .ip2(\cache_data_B[4][75] ), .op(n10833) );
  nand3_1 U13696 ( .ip1(n10835), .ip2(n10834), .ip3(n10833), .op(n12800) );
  nand2_1 U13697 ( .ip1(n12580), .ip2(n12800), .op(n10866) );
  nand2_1 U13698 ( .ip1(\cache_data_B[0][43] ), .ip2(n12204), .op(n10844) );
  and2_1 U13699 ( .ip1(n12591), .ip2(\cache_data_B[3][43] ), .op(n10841) );
  nand2_1 U13700 ( .ip1(n12584), .ip2(\cache_data_B[4][43] ), .op(n10839) );
  nand2_1 U13701 ( .ip1(n11311), .ip2(\cache_data_B[1][43] ), .op(n10838) );
  nand2_1 U13702 ( .ip1(n11296), .ip2(\cache_data_B[5][43] ), .op(n10837) );
  nand2_1 U13703 ( .ip1(n10575), .ip2(\cache_data_B[7][43] ), .op(n10836) );
  nand4_1 U13704 ( .ip1(n10839), .ip2(n10838), .ip3(n10837), .ip4(n10836), 
        .op(n10840) );
  not_ab_or_c_or_d U13705 ( .ip1(n12551), .ip2(\cache_data_B[6][43] ), .ip3(
        n10841), .ip4(n10840), .op(n10843) );
  nand2_1 U13706 ( .ip1(n11142), .ip2(\cache_data_B[2][43] ), .op(n10842) );
  nand3_1 U13707 ( .ip1(n10844), .ip2(n10843), .ip3(n10842), .op(n12812) );
  nand2_1 U13708 ( .ip1(n12563), .ip2(n12812), .op(n10865) );
  nand2_1 U13709 ( .ip1(n12559), .ip2(\cache_data_B[3][11] ), .op(n10853) );
  and2_1 U13710 ( .ip1(n12486), .ip2(\cache_data_B[2][11] ), .op(n10850) );
  nand2_1 U13711 ( .ip1(n12320), .ip2(\cache_data_B[6][11] ), .op(n10848) );
  nand2_1 U13712 ( .ip1(n12584), .ip2(\cache_data_B[4][11] ), .op(n10847) );
  nand2_1 U13713 ( .ip1(n11057), .ip2(\cache_data_B[7][11] ), .op(n10846) );
  nand2_1 U13714 ( .ip1(n11236), .ip2(\cache_data_B[5][11] ), .op(n10845) );
  nand4_1 U13715 ( .ip1(n10848), .ip2(n10847), .ip3(n10846), .ip4(n10845), 
        .op(n10849) );
  not_ab_or_c_or_d U13716 ( .ip1(\cache_data_B[0][11] ), .ip2(n8452), .ip3(
        n10850), .ip4(n10849), .op(n10852) );
  nand2_1 U13717 ( .ip1(n11311), .ip2(\cache_data_B[1][11] ), .op(n10851) );
  nand3_1 U13718 ( .ip1(n10853), .ip2(n10852), .ip3(n10851), .op(n12804) );
  nand2_1 U13719 ( .ip1(n12539), .ip2(n12804), .op(n10864) );
  nand2_1 U13720 ( .ip1(n11142), .ip2(\cache_data_B[2][107] ), .op(n10862) );
  and2_1 U13721 ( .ip1(n11946), .ip2(\cache_data_B[1][107] ), .op(n10859) );
  nand2_1 U13722 ( .ip1(n12357), .ip2(\cache_data_B[0][107] ), .op(n10857) );
  nand2_1 U13723 ( .ip1(n10702), .ip2(\cache_data_B[7][107] ), .op(n10856) );
  nand2_1 U13724 ( .ip1(n11535), .ip2(\cache_data_B[3][107] ), .op(n10855) );
  nand2_1 U13725 ( .ip1(n11236), .ip2(\cache_data_B[5][107] ), .op(n10854) );
  nand4_1 U13726 ( .ip1(n10857), .ip2(n10856), .ip3(n10855), .ip4(n10854), 
        .op(n10858) );
  not_ab_or_c_or_d U13727 ( .ip1(\cache_data_B[4][107] ), .ip2(n12476), .ip3(
        n10859), .ip4(n10858), .op(n10861) );
  nand2_1 U13728 ( .ip1(n12337), .ip2(\cache_data_B[6][107] ), .op(n10860) );
  nand3_1 U13729 ( .ip1(n10862), .ip2(n10861), .ip3(n10860), .op(n12813) );
  nand2_1 U13730 ( .ip1(n12573), .ip2(n12813), .op(n10863) );
  nand4_1 U13731 ( .ip1(n10866), .ip2(n10865), .ip3(n10864), .ip4(n10863), 
        .op(n10867) );
  not_ab_or_c_or_d U13732 ( .ip1(n12550), .ip2(n12803), .ip3(n10868), .ip4(
        n10867), .op(n10879) );
  nand2_1 U13733 ( .ip1(\cache_data_A[4][43] ), .ip2(n12584), .op(n10877) );
  and2_1 U13734 ( .ip1(n12468), .ip2(\cache_data_A[7][43] ), .op(n10874) );
  nand2_1 U13735 ( .ip1(n12320), .ip2(\cache_data_A[6][43] ), .op(n10872) );
  nand2_1 U13736 ( .ip1(n12357), .ip2(\cache_data_A[0][43] ), .op(n10871) );
  nand2_1 U13737 ( .ip1(n11296), .ip2(\cache_data_A[5][43] ), .op(n10870) );
  nand2_1 U13738 ( .ip1(n12096), .ip2(\cache_data_A[3][43] ), .op(n10869) );
  nand4_1 U13739 ( .ip1(n10872), .ip2(n10871), .ip3(n10870), .ip4(n10869), 
        .op(n10873) );
  not_ab_or_c_or_d U13740 ( .ip1(n12546), .ip2(\cache_data_A[2][43] ), .ip3(
        n10874), .ip4(n10873), .op(n10876) );
  nand2_1 U13741 ( .ip1(n11311), .ip2(\cache_data_A[1][43] ), .op(n10875) );
  nand3_1 U13742 ( .ip1(n10877), .ip2(n10876), .ip3(n10875), .op(n12802) );
  nand2_1 U13743 ( .ip1(n12595), .ip2(n12802), .op(n10878) );
  nand3_1 U13744 ( .ip1(n10880), .ip2(n10879), .ip3(n10878), .op(n10881) );
  mux2_1 U13745 ( .ip1(N4171), .ip2(n10881), .s(n11472), .op(n5309) );
  nand2_1 U13746 ( .ip1(\cache_data_B[3][108] ), .ip2(n12410), .op(n10890) );
  and2_1 U13747 ( .ip1(n12458), .ip2(\cache_data_B[6][108] ), .op(n10887) );
  nand2_1 U13748 ( .ip1(n12468), .ip2(\cache_data_B[7][108] ), .op(n10885) );
  nand2_1 U13749 ( .ip1(n11324), .ip2(\cache_data_B[4][108] ), .op(n10884) );
  nand2_1 U13750 ( .ip1(n11142), .ip2(\cache_data_B[2][108] ), .op(n10883) );
  nand2_1 U13751 ( .ip1(n11311), .ip2(\cache_data_B[1][108] ), .op(n10882) );
  nand4_1 U13752 ( .ip1(n10885), .ip2(n10884), .ip3(n10883), .ip4(n10882), 
        .op(n10886) );
  not_ab_or_c_or_d U13753 ( .ip1(\cache_data_B[0][108] ), .ip2(n12204), .ip3(
        n10887), .ip4(n10886), .op(n10889) );
  nand2_1 U13754 ( .ip1(n11296), .ip2(\cache_data_B[5][108] ), .op(n10888) );
  nand3_1 U13755 ( .ip1(n10890), .ip2(n10889), .ip3(n10888), .op(n12818) );
  nand2_1 U13756 ( .ip1(n12573), .ip2(n12818), .op(n10963) );
  nand2_1 U13757 ( .ip1(n12357), .ip2(\cache_data_B[0][44] ), .op(n10899) );
  and2_1 U13758 ( .ip1(n11946), .ip2(\cache_data_B[1][44] ), .op(n10896) );
  nand2_1 U13759 ( .ip1(n12584), .ip2(\cache_data_B[4][44] ), .op(n10894) );
  nand2_1 U13760 ( .ip1(n12320), .ip2(\cache_data_B[6][44] ), .op(n10893) );
  nand2_1 U13761 ( .ip1(n11535), .ip2(\cache_data_B[3][44] ), .op(n10892) );
  nand2_1 U13762 ( .ip1(n11296), .ip2(\cache_data_B[5][44] ), .op(n10891) );
  nand4_1 U13763 ( .ip1(n10894), .ip2(n10893), .ip3(n10892), .ip4(n10891), 
        .op(n10895) );
  not_ab_or_c_or_d U13764 ( .ip1(\cache_data_B[2][44] ), .ip2(n12546), .ip3(
        n10896), .ip4(n10895), .op(n10898) );
  nand2_1 U13765 ( .ip1(n12552), .ip2(\cache_data_B[7][44] ), .op(n10897) );
  nand3_1 U13766 ( .ip1(n10899), .ip2(n10898), .ip3(n10897), .op(n12821) );
  nand2_1 U13767 ( .ip1(n12468), .ip2(\cache_data_A[7][76] ), .op(n10903) );
  nand2_1 U13768 ( .ip1(n12096), .ip2(\cache_data_A[3][76] ), .op(n10902) );
  nand2_1 U13769 ( .ip1(n12054), .ip2(\cache_data_A[4][76] ), .op(n10901) );
  nand2_1 U13770 ( .ip1(n11311), .ip2(\cache_data_A[1][76] ), .op(n10900) );
  nand4_1 U13771 ( .ip1(n10903), .ip2(n10902), .ip3(n10901), .ip4(n10900), 
        .op(n10909) );
  nand2_1 U13772 ( .ip1(n11236), .ip2(\cache_data_A[5][76] ), .op(n10907) );
  nand2_1 U13773 ( .ip1(n11780), .ip2(\cache_data_A[6][76] ), .op(n10906) );
  nand2_1 U13774 ( .ip1(n11142), .ip2(\cache_data_A[2][76] ), .op(n10905) );
  nand2_1 U13775 ( .ip1(n12357), .ip2(\cache_data_A[0][76] ), .op(n10904) );
  nand4_1 U13776 ( .ip1(n10907), .ip2(n10906), .ip3(n10905), .ip4(n10904), 
        .op(n10908) );
  nor2_1 U13777 ( .ip1(n10909), .ip2(n10908), .op(n12819) );
  nor2_1 U13778 ( .ip1(n12819), .ip2(n12529), .op(n10951) );
  nand2_1 U13779 ( .ip1(n12357), .ip2(\cache_data_B[0][76] ), .op(n10918) );
  and2_1 U13780 ( .ip1(n12256), .ip2(\cache_data_B[5][76] ), .op(n10915) );
  nand2_1 U13781 ( .ip1(n11780), .ip2(\cache_data_B[6][76] ), .op(n10913) );
  nand2_1 U13782 ( .ip1(n12584), .ip2(\cache_data_B[4][76] ), .op(n10912) );
  nand2_1 U13783 ( .ip1(n11311), .ip2(\cache_data_B[1][76] ), .op(n10911) );
  nand2_1 U13784 ( .ip1(n12096), .ip2(\cache_data_B[3][76] ), .op(n10910) );
  nand4_1 U13785 ( .ip1(n10913), .ip2(n10912), .ip3(n10911), .ip4(n10910), 
        .op(n10914) );
  not_ab_or_c_or_d U13786 ( .ip1(\cache_data_B[2][76] ), .ip2(n12546), .ip3(
        n10915), .ip4(n10914), .op(n10917) );
  nand2_1 U13787 ( .ip1(n12552), .ip2(\cache_data_B[7][76] ), .op(n10916) );
  nand3_1 U13788 ( .ip1(n10918), .ip2(n10917), .ip3(n10916), .op(n12820) );
  nand2_1 U13789 ( .ip1(n12580), .ip2(n12820), .op(n10949) );
  nand2_1 U13790 ( .ip1(n12559), .ip2(\cache_data_A[3][12] ), .op(n10927) );
  and2_1 U13791 ( .ip1(n12396), .ip2(\cache_data_A[4][12] ), .op(n10924) );
  nand2_1 U13792 ( .ip1(n11142), .ip2(\cache_data_A[2][12] ), .op(n10922) );
  nand2_1 U13793 ( .ip1(n12357), .ip2(\cache_data_A[0][12] ), .op(n10921) );
  nand2_1 U13794 ( .ip1(n11280), .ip2(\cache_data_A[5][12] ), .op(n10920) );
  nand2_1 U13795 ( .ip1(n12581), .ip2(\cache_data_A[7][12] ), .op(n10919) );
  nand4_1 U13796 ( .ip1(n10922), .ip2(n10921), .ip3(n10920), .ip4(n10919), 
        .op(n10923) );
  not_ab_or_c_or_d U13797 ( .ip1(\cache_data_A[6][12] ), .ip2(n12551), .ip3(
        n10924), .ip4(n10923), .op(n10926) );
  nand2_1 U13798 ( .ip1(n11311), .ip2(\cache_data_A[1][12] ), .op(n10925) );
  nand3_1 U13799 ( .ip1(n10927), .ip2(n10926), .ip3(n10925), .op(n12830) );
  nand2_1 U13800 ( .ip1(n12550), .ip2(n12830), .op(n10948) );
  nand2_1 U13801 ( .ip1(\cache_data_B[2][12] ), .ip2(n12486), .op(n10936) );
  and2_1 U13802 ( .ip1(n12256), .ip2(\cache_data_B[5][12] ), .op(n10933) );
  nand2_1 U13803 ( .ip1(n11311), .ip2(\cache_data_B[1][12] ), .op(n10931) );
  nand2_1 U13804 ( .ip1(n12357), .ip2(\cache_data_B[0][12] ), .op(n10930) );
  nand2_1 U13805 ( .ip1(n11780), .ip2(\cache_data_B[6][12] ), .op(n10929) );
  nand2_1 U13806 ( .ip1(n10702), .ip2(\cache_data_B[7][12] ), .op(n10928) );
  nand4_1 U13807 ( .ip1(n10931), .ip2(n10930), .ip3(n10929), .ip4(n10928), 
        .op(n10932) );
  not_ab_or_c_or_d U13808 ( .ip1(\cache_data_B[4][12] ), .ip2(n11156), .ip3(
        n10933), .ip4(n10932), .op(n10935) );
  nand2_1 U13809 ( .ip1(n12096), .ip2(\cache_data_B[3][12] ), .op(n10934) );
  nand3_1 U13810 ( .ip1(n10936), .ip2(n10935), .ip3(n10934), .op(n12823) );
  nand2_1 U13811 ( .ip1(n12539), .ip2(n12823), .op(n10947) );
  nand2_1 U13812 ( .ip1(n12552), .ip2(\cache_data_A[7][108] ), .op(n10945) );
  and2_1 U13813 ( .ip1(n12118), .ip2(\cache_data_A[5][108] ), .op(n10942) );
  nand2_1 U13814 ( .ip1(n12357), .ip2(\cache_data_A[0][108] ), .op(n10940) );
  nand2_1 U13815 ( .ip1(n12584), .ip2(\cache_data_A[4][108] ), .op(n10939) );
  nand2_1 U13816 ( .ip1(n11142), .ip2(\cache_data_A[2][108] ), .op(n10938) );
  nand2_1 U13817 ( .ip1(n11780), .ip2(\cache_data_A[6][108] ), .op(n10937) );
  nand4_1 U13818 ( .ip1(n10940), .ip2(n10939), .ip3(n10938), .ip4(n10937), 
        .op(n10941) );
  not_ab_or_c_or_d U13819 ( .ip1(\cache_data_A[3][108] ), .ip2(n11535), .ip3(
        n10942), .ip4(n10941), .op(n10944) );
  nand2_1 U13820 ( .ip1(n11311), .ip2(\cache_data_A[1][108] ), .op(n10943) );
  nand3_1 U13821 ( .ip1(n10945), .ip2(n10944), .ip3(n10943), .op(n12822) );
  nand2_1 U13822 ( .ip1(n12509), .ip2(n12822), .op(n10946) );
  nand4_1 U13823 ( .ip1(n10949), .ip2(n10948), .ip3(n10947), .ip4(n10946), 
        .op(n10950) );
  not_ab_or_c_or_d U13824 ( .ip1(n12563), .ip2(n12821), .ip3(n10951), .ip4(
        n10950), .op(n10962) );
  nand2_1 U13825 ( .ip1(\cache_data_A[0][44] ), .ip2(n12204), .op(n10960) );
  and2_1 U13826 ( .ip1(n12147), .ip2(\cache_data_A[1][44] ), .op(n10957) );
  nand2_1 U13827 ( .ip1(n12337), .ip2(\cache_data_A[6][44] ), .op(n10955) );
  nand2_1 U13828 ( .ip1(n11280), .ip2(\cache_data_A[5][44] ), .op(n10954) );
  nand2_1 U13829 ( .ip1(n12278), .ip2(\cache_data_A[7][44] ), .op(n10953) );
  nand2_1 U13830 ( .ip1(n12476), .ip2(\cache_data_A[4][44] ), .op(n10952) );
  nand4_1 U13831 ( .ip1(n10955), .ip2(n10954), .ip3(n10953), .ip4(n10952), 
        .op(n10956) );
  not_ab_or_c_or_d U13832 ( .ip1(\cache_data_A[3][44] ), .ip2(n12096), .ip3(
        n10957), .ip4(n10956), .op(n10959) );
  nand2_1 U13833 ( .ip1(n11142), .ip2(\cache_data_A[2][44] ), .op(n10958) );
  nand3_1 U13834 ( .ip1(n10960), .ip2(n10959), .ip3(n10958), .op(n12831) );
  nand2_1 U13835 ( .ip1(n12595), .ip2(n12831), .op(n10961) );
  nand3_1 U13836 ( .ip1(n10963), .ip2(n10962), .ip3(n10961), .op(n10964) );
  mux2_1 U13837 ( .ip1(N4168), .ip2(n10964), .s(n11472), .op(n5308) );
  nand2_1 U13838 ( .ip1(n12468), .ip2(\cache_data_B[7][45] ), .op(n10973) );
  and2_1 U13839 ( .ip1(n12476), .ip2(\cache_data_B[4][45] ), .op(n10970) );
  nand2_1 U13840 ( .ip1(n11142), .ip2(\cache_data_B[2][45] ), .op(n10968) );
  nand2_1 U13841 ( .ip1(n11311), .ip2(\cache_data_B[1][45] ), .op(n10967) );
  nand2_1 U13842 ( .ip1(n12357), .ip2(\cache_data_B[0][45] ), .op(n10966) );
  nand2_1 U13843 ( .ip1(n12320), .ip2(\cache_data_B[6][45] ), .op(n10965) );
  nand4_1 U13844 ( .ip1(n10968), .ip2(n10967), .ip3(n10966), .ip4(n10965), 
        .op(n10969) );
  not_ab_or_c_or_d U13845 ( .ip1(\cache_data_B[3][45] ), .ip2(n12096), .ip3(
        n10970), .ip4(n10969), .op(n10972) );
  nand2_1 U13846 ( .ip1(n11280), .ip2(\cache_data_B[5][45] ), .op(n10971) );
  nand3_1 U13847 ( .ip1(n10973), .ip2(n10972), .ip3(n10971), .op(n12841) );
  nand2_1 U13848 ( .ip1(n12563), .ip2(n12841), .op(n11046) );
  nand2_1 U13849 ( .ip1(n12357), .ip2(\cache_data_B[0][109] ), .op(n10982) );
  and2_1 U13850 ( .ip1(n12396), .ip2(\cache_data_B[4][109] ), .op(n10979) );
  nand2_1 U13851 ( .ip1(n12096), .ip2(\cache_data_B[3][109] ), .op(n10977) );
  nand2_1 U13852 ( .ip1(n11296), .ip2(\cache_data_B[5][109] ), .op(n10976) );
  nand2_1 U13853 ( .ip1(n11142), .ip2(\cache_data_B[2][109] ), .op(n10975) );
  nand2_1 U13854 ( .ip1(n12278), .ip2(\cache_data_B[7][109] ), .op(n10974) );
  nand4_1 U13855 ( .ip1(n10977), .ip2(n10976), .ip3(n10975), .ip4(n10974), 
        .op(n10978) );
  not_ab_or_c_or_d U13856 ( .ip1(\cache_data_B[6][109] ), .ip2(n12320), .ip3(
        n10979), .ip4(n10978), .op(n10981) );
  nand2_1 U13857 ( .ip1(n11311), .ip2(\cache_data_B[1][109] ), .op(n10980) );
  nand3_1 U13858 ( .ip1(n10982), .ip2(n10981), .ip3(n10980), .op(n12849) );
  nand2_1 U13859 ( .ip1(n11142), .ip2(\cache_data_A[2][77] ), .op(n10986) );
  nand2_1 U13860 ( .ip1(n12357), .ip2(\cache_data_A[0][77] ), .op(n10985) );
  nand2_1 U13861 ( .ip1(n11236), .ip2(\cache_data_A[5][77] ), .op(n10984) );
  nand2_1 U13862 ( .ip1(n12559), .ip2(\cache_data_A[3][77] ), .op(n10983) );
  nand4_1 U13863 ( .ip1(n10986), .ip2(n10985), .ip3(n10984), .ip4(n10983), 
        .op(n10992) );
  nand2_1 U13864 ( .ip1(n12551), .ip2(\cache_data_A[6][77] ), .op(n10990) );
  nand2_1 U13865 ( .ip1(n11311), .ip2(\cache_data_A[1][77] ), .op(n10989) );
  nand2_1 U13866 ( .ip1(n11324), .ip2(\cache_data_A[4][77] ), .op(n10988) );
  nand2_1 U13867 ( .ip1(n12278), .ip2(\cache_data_A[7][77] ), .op(n10987) );
  nand4_1 U13868 ( .ip1(n10990), .ip2(n10989), .ip3(n10988), .ip4(n10987), 
        .op(n10991) );
  nor2_1 U13869 ( .ip1(n10992), .ip2(n10991), .op(n12837) );
  nor2_1 U13870 ( .ip1(n12837), .ip2(n12529), .op(n11034) );
  nand2_1 U13871 ( .ip1(n11311), .ip2(\cache_data_B[1][77] ), .op(n11001) );
  and2_1 U13872 ( .ip1(n12591), .ip2(\cache_data_B[3][77] ), .op(n10998) );
  nand2_1 U13873 ( .ip1(n12337), .ip2(\cache_data_B[6][77] ), .op(n10996) );
  nand2_1 U13874 ( .ip1(n11057), .ip2(\cache_data_B[7][77] ), .op(n10995) );
  nand2_1 U13875 ( .ip1(n11156), .ip2(\cache_data_B[4][77] ), .op(n10994) );
  nand2_1 U13876 ( .ip1(n11142), .ip2(\cache_data_B[2][77] ), .op(n10993) );
  nand4_1 U13877 ( .ip1(n10996), .ip2(n10995), .ip3(n10994), .ip4(n10993), 
        .op(n10997) );
  not_ab_or_c_or_d U13878 ( .ip1(n12297), .ip2(\cache_data_B[0][77] ), .ip3(
        n10998), .ip4(n10997), .op(n11000) );
  nand2_1 U13879 ( .ip1(n11236), .ip2(\cache_data_B[5][77] ), .op(n10999) );
  nand3_1 U13880 ( .ip1(n11001), .ip2(n11000), .ip3(n10999), .op(n12840) );
  nand2_1 U13881 ( .ip1(n12580), .ip2(n12840), .op(n11032) );
  nand2_1 U13882 ( .ip1(n12551), .ip2(\cache_data_A[6][109] ), .op(n11010) );
  and2_1 U13883 ( .ip1(n12321), .ip2(\cache_data_A[3][109] ), .op(n11007) );
  nand2_1 U13884 ( .ip1(n11311), .ip2(\cache_data_A[1][109] ), .op(n11005) );
  nand2_1 U13885 ( .ip1(n11156), .ip2(\cache_data_A[4][109] ), .op(n11004) );
  nand2_1 U13886 ( .ip1(n12468), .ip2(\cache_data_A[7][109] ), .op(n11003) );
  nand2_1 U13887 ( .ip1(n12357), .ip2(\cache_data_A[0][109] ), .op(n11002) );
  nand4_1 U13888 ( .ip1(n11005), .ip2(n11004), .ip3(n11003), .ip4(n11002), 
        .op(n11006) );
  not_ab_or_c_or_d U13889 ( .ip1(\cache_data_A[2][109] ), .ip2(n12475), .ip3(
        n11007), .ip4(n11006), .op(n11009) );
  nand2_1 U13890 ( .ip1(n11304), .ip2(\cache_data_A[5][109] ), .op(n11008) );
  nand3_1 U13891 ( .ip1(n11010), .ip2(n11009), .ip3(n11008), .op(n12838) );
  nand2_1 U13892 ( .ip1(n12509), .ip2(n12838), .op(n11031) );
  nand2_1 U13893 ( .ip1(n12559), .ip2(\cache_data_A[3][13] ), .op(n11019) );
  and2_1 U13894 ( .ip1(n12581), .ip2(\cache_data_A[7][13] ), .op(n11016) );
  nand2_1 U13895 ( .ip1(n11142), .ip2(\cache_data_A[2][13] ), .op(n11014) );
  nand2_1 U13896 ( .ip1(n11156), .ip2(\cache_data_A[4][13] ), .op(n11013) );
  nand2_1 U13897 ( .ip1(n11311), .ip2(\cache_data_A[1][13] ), .op(n11012) );
  nand2_1 U13898 ( .ip1(n12337), .ip2(\cache_data_A[6][13] ), .op(n11011) );
  nand4_1 U13899 ( .ip1(n11014), .ip2(n11013), .ip3(n11012), .ip4(n11011), 
        .op(n11015) );
  not_ab_or_c_or_d U13900 ( .ip1(n12297), .ip2(\cache_data_A[0][13] ), .ip3(
        n11016), .ip4(n11015), .op(n11018) );
  nand2_1 U13901 ( .ip1(n11280), .ip2(\cache_data_A[5][13] ), .op(n11017) );
  nand3_1 U13902 ( .ip1(n11019), .ip2(n11018), .ip3(n11017), .op(n12848) );
  nand2_1 U13903 ( .ip1(n12550), .ip2(n12848), .op(n11030) );
  nand2_1 U13904 ( .ip1(\cache_data_A[7][45] ), .ip2(n12468), .op(n11028) );
  and2_1 U13905 ( .ip1(n12486), .ip2(\cache_data_A[2][45] ), .op(n11025) );
  nand2_1 U13906 ( .ip1(n12096), .ip2(\cache_data_A[3][45] ), .op(n11023) );
  nand2_1 U13907 ( .ip1(n11311), .ip2(\cache_data_A[1][45] ), .op(n11022) );
  nand2_1 U13908 ( .ip1(n12054), .ip2(\cache_data_A[4][45] ), .op(n11021) );
  nand2_1 U13909 ( .ip1(n12337), .ip2(\cache_data_A[6][45] ), .op(n11020) );
  nand4_1 U13910 ( .ip1(n11023), .ip2(n11022), .ip3(n11021), .ip4(n11020), 
        .op(n11024) );
  not_ab_or_c_or_d U13911 ( .ip1(\cache_data_A[0][45] ), .ip2(n12357), .ip3(
        n11025), .ip4(n11024), .op(n11027) );
  nand2_1 U13912 ( .ip1(n11280), .ip2(\cache_data_A[5][45] ), .op(n11026) );
  nand3_1 U13913 ( .ip1(n11028), .ip2(n11027), .ip3(n11026), .op(n12836) );
  nand2_1 U13914 ( .ip1(n12595), .ip2(n12836), .op(n11029) );
  nand4_1 U13915 ( .ip1(n11032), .ip2(n11031), .ip3(n11030), .ip4(n11029), 
        .op(n11033) );
  not_ab_or_c_or_d U13916 ( .ip1(n12573), .ip2(n12849), .ip3(n11034), .ip4(
        n11033), .op(n11045) );
  nand2_1 U13917 ( .ip1(n11324), .ip2(\cache_data_B[4][13] ), .op(n11043) );
  and2_1 U13918 ( .ip1(n8060), .ip2(\cache_data_B[3][13] ), .op(n11040) );
  nand2_1 U13919 ( .ip1(n12320), .ip2(\cache_data_B[6][13] ), .op(n11038) );
  nand2_1 U13920 ( .ip1(n11142), .ip2(\cache_data_B[2][13] ), .op(n11037) );
  nand2_1 U13921 ( .ip1(n11057), .ip2(\cache_data_B[7][13] ), .op(n11036) );
  nand2_1 U13922 ( .ip1(n11304), .ip2(\cache_data_B[5][13] ), .op(n11035) );
  nand4_1 U13923 ( .ip1(n11038), .ip2(n11037), .ip3(n11036), .ip4(n11035), 
        .op(n11039) );
  not_ab_or_c_or_d U13924 ( .ip1(\cache_data_B[0][13] ), .ip2(n12357), .ip3(
        n11040), .ip4(n11039), .op(n11042) );
  nand2_1 U13925 ( .ip1(n11311), .ip2(\cache_data_B[1][13] ), .op(n11041) );
  nand3_1 U13926 ( .ip1(n11043), .ip2(n11042), .ip3(n11041), .op(n12839) );
  nand2_1 U13927 ( .ip1(n12539), .ip2(n12839), .op(n11044) );
  nand3_1 U13928 ( .ip1(n11046), .ip2(n11045), .ip3(n11044), .op(n11047) );
  mux2_1 U13929 ( .ip1(N4165), .ip2(n11047), .s(n11472), .op(n5307) );
  nand2_1 U13930 ( .ip1(n12458), .ip2(\cache_data_B[6][110] ), .op(n11056) );
  and2_1 U13931 ( .ip1(n12581), .ip2(\cache_data_B[7][110] ), .op(n11053) );
  nand2_1 U13932 ( .ip1(n11142), .ip2(\cache_data_B[2][110] ), .op(n11051) );
  nand2_1 U13933 ( .ip1(n12559), .ip2(\cache_data_B[3][110] ), .op(n11050) );
  nand2_1 U13934 ( .ip1(n11311), .ip2(\cache_data_B[1][110] ), .op(n11049) );
  nand2_1 U13935 ( .ip1(n11324), .ip2(\cache_data_B[4][110] ), .op(n11048) );
  nand4_1 U13936 ( .ip1(n11051), .ip2(n11050), .ip3(n11049), .ip4(n11048), 
        .op(n11052) );
  not_ab_or_c_or_d U13937 ( .ip1(\cache_data_B[0][110] ), .ip2(n12204), .ip3(
        n11053), .ip4(n11052), .op(n11055) );
  nand2_1 U13938 ( .ip1(n11236), .ip2(\cache_data_B[5][110] ), .op(n11054) );
  nand3_1 U13939 ( .ip1(n11056), .ip2(n11055), .ip3(n11054), .op(n12866) );
  nand2_1 U13940 ( .ip1(n12573), .ip2(n12866), .op(n11131) );
  nand2_1 U13941 ( .ip1(\cache_data_A[0][14] ), .ip2(n12204), .op(n11066) );
  and2_1 U13942 ( .ip1(n12582), .ip2(\cache_data_A[5][14] ), .op(n11063) );
  nand2_1 U13943 ( .ip1(n12584), .ip2(\cache_data_A[4][14] ), .op(n11061) );
  nand2_1 U13944 ( .ip1(n11311), .ip2(\cache_data_A[1][14] ), .op(n11060) );
  nand2_1 U13945 ( .ip1(n11057), .ip2(\cache_data_A[7][14] ), .op(n11059) );
  nand2_1 U13946 ( .ip1(n12458), .ip2(\cache_data_A[6][14] ), .op(n11058) );
  nand4_1 U13947 ( .ip1(n11061), .ip2(n11060), .ip3(n11059), .ip4(n11058), 
        .op(n11062) );
  not_ab_or_c_or_d U13948 ( .ip1(\cache_data_A[2][14] ), .ip2(n12546), .ip3(
        n11063), .ip4(n11062), .op(n11065) );
  nand2_1 U13949 ( .ip1(n12096), .ip2(\cache_data_A[3][14] ), .op(n11064) );
  nand3_1 U13950 ( .ip1(n11066), .ip2(n11065), .ip3(n11064), .op(n12856) );
  nand2_1 U13951 ( .ip1(n12278), .ip2(\cache_data_A[7][78] ), .op(n11070) );
  nand2_1 U13952 ( .ip1(n11311), .ip2(\cache_data_A[1][78] ), .op(n11069) );
  nand2_1 U13953 ( .ip1(n12551), .ip2(\cache_data_A[6][78] ), .op(n11068) );
  nand2_1 U13954 ( .ip1(n12559), .ip2(\cache_data_A[3][78] ), .op(n11067) );
  nand4_1 U13955 ( .ip1(n11070), .ip2(n11069), .ip3(n11068), .ip4(n11067), 
        .op(n11077) );
  nand2_1 U13956 ( .ip1(n11156), .ip2(\cache_data_A[4][78] ), .op(n11075) );
  nand2_1 U13957 ( .ip1(n12546), .ip2(\cache_data_A[2][78] ), .op(n11074) );
  nand2_1 U13958 ( .ip1(n11071), .ip2(\cache_data_A[0][78] ), .op(n11073) );
  nand2_1 U13959 ( .ip1(n11280), .ip2(\cache_data_A[5][78] ), .op(n11072) );
  nand4_1 U13960 ( .ip1(n11075), .ip2(n11074), .ip3(n11073), .ip4(n11072), 
        .op(n11076) );
  nor2_1 U13961 ( .ip1(n11077), .ip2(n11076), .op(n12855) );
  nor2_1 U13962 ( .ip1(n12855), .ip2(n12529), .op(n11119) );
  nand2_1 U13963 ( .ip1(n12468), .ip2(\cache_data_B[7][14] ), .op(n11086) );
  and2_1 U13964 ( .ip1(n12429), .ip2(\cache_data_B[6][14] ), .op(n11083) );
  nand2_1 U13965 ( .ip1(n11535), .ip2(\cache_data_B[3][14] ), .op(n11081) );
  nand2_1 U13966 ( .ip1(n11311), .ip2(\cache_data_B[1][14] ), .op(n11080) );
  nand2_1 U13967 ( .ip1(n12475), .ip2(\cache_data_B[2][14] ), .op(n11079) );
  nand2_1 U13968 ( .ip1(n12584), .ip2(\cache_data_B[4][14] ), .op(n11078) );
  nand4_1 U13969 ( .ip1(n11081), .ip2(n11080), .ip3(n11079), .ip4(n11078), 
        .op(n11082) );
  not_ab_or_c_or_d U13970 ( .ip1(\cache_data_B[0][14] ), .ip2(n11911), .ip3(
        n11083), .ip4(n11082), .op(n11085) );
  nand2_1 U13971 ( .ip1(n11304), .ip2(\cache_data_B[5][14] ), .op(n11084) );
  nand3_1 U13972 ( .ip1(n11086), .ip2(n11085), .ip3(n11084), .op(n12858) );
  nand2_1 U13973 ( .ip1(n12539), .ip2(n12858), .op(n11117) );
  nand2_1 U13974 ( .ip1(n12337), .ip2(\cache_data_B[6][78] ), .op(n11095) );
  and2_1 U13975 ( .ip1(n12321), .ip2(\cache_data_B[3][78] ), .op(n11092) );
  nand2_1 U13976 ( .ip1(n11304), .ip2(\cache_data_B[5][78] ), .op(n11090) );
  nand2_1 U13977 ( .ip1(n11142), .ip2(\cache_data_B[2][78] ), .op(n11089) );
  nand2_1 U13978 ( .ip1(n12054), .ip2(\cache_data_B[4][78] ), .op(n11088) );
  nand2_1 U13979 ( .ip1(n10702), .ip2(\cache_data_B[7][78] ), .op(n11087) );
  nand4_1 U13980 ( .ip1(n11090), .ip2(n11089), .ip3(n11088), .ip4(n11087), 
        .op(n11091) );
  not_ab_or_c_or_d U13981 ( .ip1(\cache_data_B[0][78] ), .ip2(n12357), .ip3(
        n11092), .ip4(n11091), .op(n11094) );
  nand2_1 U13982 ( .ip1(n11311), .ip2(\cache_data_B[1][78] ), .op(n11093) );
  nand3_1 U13983 ( .ip1(n11095), .ip2(n11094), .ip3(n11093), .op(n12857) );
  nand2_1 U13984 ( .ip1(n12580), .ip2(n12857), .op(n11116) );
  nand2_1 U13985 ( .ip1(\cache_data_B[7][46] ), .ip2(n12468), .op(n11104) );
  and2_1 U13986 ( .ip1(n11946), .ip2(\cache_data_B[1][46] ), .op(n11101) );
  buf_1 U13987 ( .ip(n12370), .op(n11911) );
  nand2_1 U13988 ( .ip1(n11911), .ip2(\cache_data_B[0][46] ), .op(n11099) );
  nand2_1 U13989 ( .ip1(n11280), .ip2(\cache_data_B[5][46] ), .op(n11098) );
  nand2_1 U13990 ( .ip1(n12584), .ip2(\cache_data_B[4][46] ), .op(n11097) );
  nand2_1 U13991 ( .ip1(n12475), .ip2(\cache_data_B[2][46] ), .op(n11096) );
  nand4_1 U13992 ( .ip1(n11099), .ip2(n11098), .ip3(n11097), .ip4(n11096), 
        .op(n11100) );
  not_ab_or_c_or_d U13993 ( .ip1(n12096), .ip2(\cache_data_B[3][46] ), .ip3(
        n11101), .ip4(n11100), .op(n11103) );
  nand2_1 U13994 ( .ip1(n12551), .ip2(\cache_data_B[6][46] ), .op(n11102) );
  nand3_1 U13995 ( .ip1(n11104), .ip2(n11103), .ip3(n11102), .op(n12859) );
  nand2_1 U13996 ( .ip1(n12563), .ip2(n12859), .op(n11115) );
  nand2_1 U13997 ( .ip1(n11535), .ip2(\cache_data_A[3][110] ), .op(n11113) );
  and2_1 U13998 ( .ip1(n11946), .ip2(\cache_data_A[1][110] ), .op(n11110) );
  nand2_1 U13999 ( .ip1(n12204), .ip2(\cache_data_A[0][110] ), .op(n11108) );
  nand2_1 U14000 ( .ip1(n10702), .ip2(\cache_data_A[7][110] ), .op(n11107) );
  nand2_1 U14001 ( .ip1(n12337), .ip2(\cache_data_A[6][110] ), .op(n11106) );
  nand2_1 U14002 ( .ip1(n11304), .ip2(\cache_data_A[5][110] ), .op(n11105) );
  nand4_1 U14003 ( .ip1(n11108), .ip2(n11107), .ip3(n11106), .ip4(n11105), 
        .op(n11109) );
  not_ab_or_c_or_d U14004 ( .ip1(\cache_data_A[2][110] ), .ip2(n12475), .ip3(
        n11110), .ip4(n11109), .op(n11112) );
  nand2_1 U14005 ( .ip1(n11324), .ip2(\cache_data_A[4][110] ), .op(n11111) );
  nand3_1 U14006 ( .ip1(n11113), .ip2(n11112), .ip3(n11111), .op(n12854) );
  nand2_1 U14007 ( .ip1(n12509), .ip2(n12854), .op(n11114) );
  nand4_1 U14008 ( .ip1(n11117), .ip2(n11116), .ip3(n11115), .ip4(n11114), 
        .op(n11118) );
  not_ab_or_c_or_d U14009 ( .ip1(n12550), .ip2(n12856), .ip3(n11119), .ip4(
        n11118), .op(n11130) );
  nand2_1 U14010 ( .ip1(\cache_data_A[7][46] ), .ip2(n12552), .op(n11128) );
  and2_1 U14011 ( .ip1(n11296), .ip2(\cache_data_A[5][46] ), .op(n11125) );
  nand2_1 U14012 ( .ip1(n11324), .ip2(\cache_data_A[4][46] ), .op(n11123) );
  nand2_1 U14013 ( .ip1(n12096), .ip2(\cache_data_A[3][46] ), .op(n11122) );
  nand2_1 U14014 ( .ip1(n11311), .ip2(\cache_data_A[1][46] ), .op(n11121) );
  nand2_1 U14015 ( .ip1(n11142), .ip2(\cache_data_A[2][46] ), .op(n11120) );
  nand4_1 U14016 ( .ip1(n11123), .ip2(n11122), .ip3(n11121), .ip4(n11120), 
        .op(n11124) );
  not_ab_or_c_or_d U14017 ( .ip1(\cache_data_A[0][46] ), .ip2(n12357), .ip3(
        n11125), .ip4(n11124), .op(n11127) );
  nand2_1 U14018 ( .ip1(n12320), .ip2(\cache_data_A[6][46] ), .op(n11126) );
  nand3_1 U14019 ( .ip1(n11128), .ip2(n11127), .ip3(n11126), .op(n12867) );
  nand2_1 U14020 ( .ip1(n12595), .ip2(n12867), .op(n11129) );
  nand3_1 U14021 ( .ip1(n11131), .ip2(n11130), .ip3(n11129), .op(n11132) );
  mux2_1 U14022 ( .ip1(N4162), .ip2(n11132), .s(n11472), .op(n5306) );
  nand2_1 U14023 ( .ip1(n12552), .ip2(\cache_data_B[7][111] ), .op(n11141) );
  and2_1 U14024 ( .ip1(n12476), .ip2(\cache_data_B[4][111] ), .op(n11138) );
  nand2_1 U14025 ( .ip1(n12475), .ip2(\cache_data_B[2][111] ), .op(n11136) );
  nand2_1 U14026 ( .ip1(n11304), .ip2(\cache_data_B[5][111] ), .op(n11135) );
  nand2_1 U14027 ( .ip1(n12204), .ip2(\cache_data_B[0][111] ), .op(n11134) );
  nand2_1 U14028 ( .ip1(n11311), .ip2(\cache_data_B[1][111] ), .op(n11133) );
  nand4_1 U14029 ( .ip1(n11136), .ip2(n11135), .ip3(n11134), .ip4(n11133), 
        .op(n11137) );
  not_ab_or_c_or_d U14030 ( .ip1(n12551), .ip2(\cache_data_B[6][111] ), .ip3(
        n11138), .ip4(n11137), .op(n11140) );
  nand2_1 U14031 ( .ip1(n12096), .ip2(\cache_data_B[3][111] ), .op(n11139) );
  nand3_1 U14032 ( .ip1(n11141), .ip2(n11140), .ip3(n11139), .op(n12874) );
  nand2_1 U14033 ( .ip1(n12573), .ip2(n12874), .op(n11216) );
  nand2_1 U14034 ( .ip1(n11311), .ip2(\cache_data_A[1][111] ), .op(n11151) );
  and2_1 U14035 ( .ip1(n12458), .ip2(\cache_data_A[6][111] ), .op(n11148) );
  nand2_1 U14036 ( .ip1(n11142), .ip2(\cache_data_A[2][111] ), .op(n11146) );
  nand2_1 U14037 ( .ip1(n12054), .ip2(\cache_data_A[4][111] ), .op(n11145) );
  nand2_1 U14038 ( .ip1(n11911), .ip2(\cache_data_A[0][111] ), .op(n11144) );
  nand2_1 U14039 ( .ip1(n12559), .ip2(\cache_data_A[3][111] ), .op(n11143) );
  nand4_1 U14040 ( .ip1(n11146), .ip2(n11145), .ip3(n11144), .ip4(n11143), 
        .op(n11147) );
  not_ab_or_c_or_d U14041 ( .ip1(\cache_data_A[7][111] ), .ip2(n12278), .ip3(
        n11148), .ip4(n11147), .op(n11150) );
  nand2_1 U14042 ( .ip1(n11296), .ip2(\cache_data_A[5][111] ), .op(n11149) );
  nand3_1 U14043 ( .ip1(n11151), .ip2(n11150), .ip3(n11149), .op(n12872) );
  nand2_1 U14044 ( .ip1(n12204), .ip2(\cache_data_A[0][79] ), .op(n11155) );
  nand2_1 U14045 ( .ip1(n12096), .ip2(\cache_data_A[3][79] ), .op(n11154) );
  nand2_1 U14046 ( .ip1(n11280), .ip2(\cache_data_A[5][79] ), .op(n11153) );
  nand2_1 U14047 ( .ip1(n10575), .ip2(\cache_data_A[7][79] ), .op(n11152) );
  nand4_1 U14048 ( .ip1(n11155), .ip2(n11154), .ip3(n11153), .ip4(n11152), 
        .op(n11162) );
  nand2_1 U14049 ( .ip1(n12551), .ip2(\cache_data_A[6][79] ), .op(n11160) );
  nand2_1 U14050 ( .ip1(n11855), .ip2(\cache_data_A[2][79] ), .op(n11159) );
  nand2_1 U14051 ( .ip1(n11156), .ip2(\cache_data_A[4][79] ), .op(n11158) );
  nand2_1 U14052 ( .ip1(n11311), .ip2(\cache_data_A[1][79] ), .op(n11157) );
  nand4_1 U14053 ( .ip1(n11160), .ip2(n11159), .ip3(n11158), .ip4(n11157), 
        .op(n11161) );
  nor2_1 U14054 ( .ip1(n11162), .ip2(n11161), .op(n12873) );
  nor2_1 U14055 ( .ip1(n12873), .ip2(n12529), .op(n11204) );
  nand2_1 U14056 ( .ip1(n12486), .ip2(\cache_data_A[2][47] ), .op(n11171) );
  and2_1 U14057 ( .ip1(n11296), .ip2(\cache_data_A[5][47] ), .op(n11168) );
  nand2_1 U14058 ( .ip1(n12320), .ip2(\cache_data_A[6][47] ), .op(n11166) );
  nand2_1 U14059 ( .ip1(n11535), .ip2(\cache_data_A[3][47] ), .op(n11165) );
  nand2_1 U14060 ( .ip1(n12204), .ip2(\cache_data_A[0][47] ), .op(n11164) );
  nand2_1 U14061 ( .ip1(n11311), .ip2(\cache_data_A[1][47] ), .op(n11163) );
  nand4_1 U14062 ( .ip1(n11166), .ip2(n11165), .ip3(n11164), .ip4(n11163), 
        .op(n11167) );
  not_ab_or_c_or_d U14063 ( .ip1(n11156), .ip2(\cache_data_A[4][47] ), .ip3(
        n11168), .ip4(n11167), .op(n11170) );
  nand2_1 U14064 ( .ip1(n12552), .ip2(\cache_data_A[7][47] ), .op(n11169) );
  nand3_1 U14065 ( .ip1(n11171), .ip2(n11170), .ip3(n11169), .op(n12885) );
  nand2_1 U14066 ( .ip1(n12595), .ip2(n12885), .op(n11202) );
  nand2_1 U14067 ( .ip1(n12096), .ip2(\cache_data_A[3][15] ), .op(n11180) );
  and2_1 U14068 ( .ip1(n12147), .ip2(\cache_data_A[1][15] ), .op(n11177) );
  nand2_1 U14069 ( .ip1(n12552), .ip2(\cache_data_A[7][15] ), .op(n11175) );
  nand2_1 U14070 ( .ip1(n12486), .ip2(\cache_data_A[2][15] ), .op(n11174) );
  nand2_1 U14071 ( .ip1(n11911), .ip2(\cache_data_A[0][15] ), .op(n11173) );
  nand2_1 U14072 ( .ip1(n11156), .ip2(\cache_data_A[4][15] ), .op(n11172) );
  nand4_1 U14073 ( .ip1(n11175), .ip2(n11174), .ip3(n11173), .ip4(n11172), 
        .op(n11176) );
  not_ab_or_c_or_d U14074 ( .ip1(\cache_data_A[6][15] ), .ip2(n12551), .ip3(
        n11177), .ip4(n11176), .op(n11179) );
  nand2_1 U14075 ( .ip1(n11304), .ip2(\cache_data_A[5][15] ), .op(n11178) );
  nand3_1 U14076 ( .ip1(n11180), .ip2(n11179), .ip3(n11178), .op(n12884) );
  nand2_1 U14077 ( .ip1(n12550), .ip2(n12884), .op(n11201) );
  nand2_1 U14078 ( .ip1(\cache_data_B[3][15] ), .ip2(n8060), .op(n11189) );
  and2_1 U14079 ( .ip1(n12486), .ip2(\cache_data_B[2][15] ), .op(n11186) );
  nand2_1 U14080 ( .ip1(n10575), .ip2(\cache_data_B[7][15] ), .op(n11184) );
  nand2_1 U14081 ( .ip1(n11304), .ip2(\cache_data_B[5][15] ), .op(n11183) );
  nand2_1 U14082 ( .ip1(n12371), .ip2(\cache_data_B[6][15] ), .op(n11182) );
  nand2_1 U14083 ( .ip1(n12054), .ip2(\cache_data_B[4][15] ), .op(n11181) );
  nand4_1 U14084 ( .ip1(n11184), .ip2(n11183), .ip3(n11182), .ip4(n11181), 
        .op(n11185) );
  not_ab_or_c_or_d U14085 ( .ip1(\cache_data_B[0][15] ), .ip2(n12357), .ip3(
        n11186), .ip4(n11185), .op(n11188) );
  nand2_1 U14086 ( .ip1(n11311), .ip2(\cache_data_B[1][15] ), .op(n11187) );
  nand3_1 U14087 ( .ip1(n11189), .ip2(n11188), .ip3(n11187), .op(n12877) );
  nand2_1 U14088 ( .ip1(n12539), .ip2(n12877), .op(n11200) );
  nand2_1 U14089 ( .ip1(n11855), .ip2(\cache_data_B[2][47] ), .op(n11198) );
  and2_1 U14090 ( .ip1(n11304), .ip2(\cache_data_B[5][47] ), .op(n11195) );
  nand2_1 U14091 ( .ip1(n12096), .ip2(\cache_data_B[3][47] ), .op(n11193) );
  nand2_1 U14092 ( .ip1(n12370), .ip2(\cache_data_B[0][47] ), .op(n11192) );
  nand2_1 U14093 ( .ip1(n10702), .ip2(\cache_data_B[7][47] ), .op(n11191) );
  nand2_1 U14094 ( .ip1(n12458), .ip2(\cache_data_B[6][47] ), .op(n11190) );
  nand4_1 U14095 ( .ip1(n11193), .ip2(n11192), .ip3(n11191), .ip4(n11190), 
        .op(n11194) );
  not_ab_or_c_or_d U14096 ( .ip1(\cache_data_B[1][47] ), .ip2(n11946), .ip3(
        n11195), .ip4(n11194), .op(n11197) );
  nand2_1 U14097 ( .ip1(n11156), .ip2(\cache_data_B[4][47] ), .op(n11196) );
  nand3_1 U14098 ( .ip1(n11198), .ip2(n11197), .ip3(n11196), .op(n12875) );
  nand2_1 U14099 ( .ip1(n12563), .ip2(n12875), .op(n11199) );
  nand4_1 U14100 ( .ip1(n11202), .ip2(n11201), .ip3(n11200), .ip4(n11199), 
        .op(n11203) );
  not_ab_or_c_or_d U14101 ( .ip1(n12509), .ip2(n12872), .ip3(n11204), .ip4(
        n11203), .op(n11215) );
  nand2_1 U14102 ( .ip1(n12337), .ip2(\cache_data_B[6][79] ), .op(n11213) );
  and2_1 U14103 ( .ip1(n12476), .ip2(\cache_data_B[4][79] ), .op(n11210) );
  nand2_1 U14104 ( .ip1(n12559), .ip2(\cache_data_B[3][79] ), .op(n11208) );
  nand2_1 U14105 ( .ip1(n12486), .ip2(\cache_data_B[2][79] ), .op(n11207) );
  nand2_1 U14106 ( .ip1(n12278), .ip2(\cache_data_B[7][79] ), .op(n11206) );
  nand2_1 U14107 ( .ip1(n11311), .ip2(\cache_data_B[1][79] ), .op(n11205) );
  nand4_1 U14108 ( .ip1(n11208), .ip2(n11207), .ip3(n11206), .ip4(n11205), 
        .op(n11209) );
  not_ab_or_c_or_d U14109 ( .ip1(n12297), .ip2(\cache_data_B[0][79] ), .ip3(
        n11210), .ip4(n11209), .op(n11212) );
  nand2_1 U14110 ( .ip1(n11280), .ip2(\cache_data_B[5][79] ), .op(n11211) );
  nand3_1 U14111 ( .ip1(n11213), .ip2(n11212), .ip3(n11211), .op(n12876) );
  nand2_1 U14112 ( .ip1(n12580), .ip2(n12876), .op(n11214) );
  nand3_1 U14113 ( .ip1(n11216), .ip2(n11215), .ip3(n11214), .op(n11217) );
  mux2_1 U14114 ( .ip1(N4159), .ip2(n11217), .s(n11472), .op(n5305) );
  nand2_1 U14115 ( .ip1(n12559), .ip2(\cache_data_A[3][16] ), .op(n11226) );
  and2_1 U14116 ( .ip1(n12486), .ip2(\cache_data_A[2][16] ), .op(n11223) );
  nand2_1 U14117 ( .ip1(n11311), .ip2(\cache_data_A[1][16] ), .op(n11221) );
  nand2_1 U14118 ( .ip1(n10575), .ip2(\cache_data_A[7][16] ), .op(n11220) );
  nand2_1 U14119 ( .ip1(n12476), .ip2(\cache_data_A[4][16] ), .op(n11219) );
  nand2_1 U14120 ( .ip1(n12320), .ip2(\cache_data_A[6][16] ), .op(n11218) );
  nand4_1 U14121 ( .ip1(n11221), .ip2(n11220), .ip3(n11219), .ip4(n11218), 
        .op(n11222) );
  not_ab_or_c_or_d U14122 ( .ip1(n12204), .ip2(\cache_data_A[0][16] ), .ip3(
        n11223), .ip4(n11222), .op(n11225) );
  nand2_1 U14123 ( .ip1(n11236), .ip2(\cache_data_A[5][16] ), .op(n11224) );
  nand3_1 U14124 ( .ip1(n11226), .ip2(n11225), .ip3(n11224), .op(n12902) );
  nand2_1 U14125 ( .ip1(n12550), .ip2(n12902), .op(n11302) );
  nand2_1 U14126 ( .ip1(\cache_data_B[4][80] ), .ip2(n12194), .op(n11235) );
  and2_1 U14127 ( .ip1(n12581), .ip2(\cache_data_B[7][80] ), .op(n11232) );
  nand2_1 U14128 ( .ip1(n11535), .ip2(\cache_data_B[3][80] ), .op(n11230) );
  nand2_1 U14129 ( .ip1(n12337), .ip2(\cache_data_B[6][80] ), .op(n11229) );
  nand2_1 U14130 ( .ip1(n11280), .ip2(\cache_data_B[5][80] ), .op(n11228) );
  nand2_1 U14131 ( .ip1(n12486), .ip2(\cache_data_B[2][80] ), .op(n11227) );
  nand4_1 U14132 ( .ip1(n11230), .ip2(n11229), .ip3(n11228), .ip4(n11227), 
        .op(n11231) );
  not_ab_or_c_or_d U14133 ( .ip1(n8452), .ip2(\cache_data_B[0][80] ), .ip3(
        n11232), .ip4(n11231), .op(n11234) );
  nand2_1 U14134 ( .ip1(n11311), .ip2(\cache_data_B[1][80] ), .op(n11233) );
  nand3_1 U14135 ( .ip1(n11235), .ip2(n11234), .ip3(n11233), .op(n12890) );
  nand2_1 U14136 ( .ip1(n11911), .ip2(\cache_data_A[0][80] ), .op(n11240) );
  nand2_1 U14137 ( .ip1(n11311), .ip2(\cache_data_A[1][80] ), .op(n11239) );
  nand2_1 U14138 ( .ip1(n11236), .ip2(\cache_data_A[5][80] ), .op(n11238) );
  nand2_1 U14139 ( .ip1(n12552), .ip2(\cache_data_A[7][80] ), .op(n11237) );
  nand4_1 U14140 ( .ip1(n11240), .ip2(n11239), .ip3(n11238), .ip4(n11237), 
        .op(n11246) );
  nand2_1 U14141 ( .ip1(n12559), .ip2(\cache_data_A[3][80] ), .op(n11244) );
  nand2_1 U14142 ( .ip1(n12429), .ip2(\cache_data_A[6][80] ), .op(n11243) );
  nand2_1 U14143 ( .ip1(n11324), .ip2(\cache_data_A[4][80] ), .op(n11242) );
  nand2_1 U14144 ( .ip1(n11855), .ip2(\cache_data_A[2][80] ), .op(n11241) );
  nand4_1 U14145 ( .ip1(n11244), .ip2(n11243), .ip3(n11242), .ip4(n11241), 
        .op(n11245) );
  nor2_1 U14146 ( .ip1(n11246), .ip2(n11245), .op(n12891) );
  nor2_1 U14147 ( .ip1(n12891), .ip2(n12529), .op(n11289) );
  nand2_1 U14148 ( .ip1(\cache_data_B[2][112] ), .ip2(n12486), .op(n11255) );
  and2_1 U14149 ( .ip1(n12476), .ip2(\cache_data_B[4][112] ), .op(n11252) );
  nand2_1 U14150 ( .ip1(n12096), .ip2(\cache_data_B[3][112] ), .op(n11250) );
  nand2_1 U14151 ( .ip1(n11280), .ip2(\cache_data_B[5][112] ), .op(n11249) );
  nand2_1 U14152 ( .ip1(n10702), .ip2(\cache_data_B[7][112] ), .op(n11248) );
  nand2_1 U14153 ( .ip1(n11946), .ip2(\cache_data_B[1][112] ), .op(n11247) );
  nand4_1 U14154 ( .ip1(n11250), .ip2(n11249), .ip3(n11248), .ip4(n11247), 
        .op(n11251) );
  not_ab_or_c_or_d U14155 ( .ip1(n12297), .ip2(\cache_data_B[0][112] ), .ip3(
        n11252), .ip4(n11251), .op(n11254) );
  nand2_1 U14156 ( .ip1(n12458), .ip2(\cache_data_B[6][112] ), .op(n11253) );
  nand3_1 U14157 ( .ip1(n11255), .ip2(n11254), .ip3(n11253), .op(n12903) );
  nand2_1 U14158 ( .ip1(n12573), .ip2(n12903), .op(n11287) );
  nand2_1 U14159 ( .ip1(n12320), .ip2(\cache_data_B[6][16] ), .op(n11264) );
  and2_1 U14160 ( .ip1(n10686), .ip2(\cache_data_B[1][16] ), .op(n11261) );
  nand2_1 U14161 ( .ip1(n11855), .ip2(\cache_data_B[2][16] ), .op(n11259) );
  nand2_1 U14162 ( .ip1(n12096), .ip2(\cache_data_B[3][16] ), .op(n11258) );
  nand2_1 U14163 ( .ip1(n12584), .ip2(\cache_data_B[4][16] ), .op(n11257) );
  nand2_1 U14164 ( .ip1(n10575), .ip2(\cache_data_B[7][16] ), .op(n11256) );
  nand4_1 U14165 ( .ip1(n11259), .ip2(n11258), .ip3(n11257), .ip4(n11256), 
        .op(n11260) );
  not_ab_or_c_or_d U14166 ( .ip1(\cache_data_B[0][16] ), .ip2(n12357), .ip3(
        n11261), .ip4(n11260), .op(n11263) );
  nand2_1 U14167 ( .ip1(n11280), .ip2(\cache_data_B[5][16] ), .op(n11262) );
  nand3_1 U14168 ( .ip1(n11264), .ip2(n11263), .ip3(n11262), .op(n12892) );
  nand2_1 U14169 ( .ip1(n12539), .ip2(n12892), .op(n11286) );
  nand2_1 U14170 ( .ip1(n11324), .ip2(\cache_data_B[4][48] ), .op(n11273) );
  and2_1 U14171 ( .ip1(n12410), .ip2(\cache_data_B[3][48] ), .op(n11270) );
  nand2_1 U14172 ( .ip1(n11311), .ip2(\cache_data_B[1][48] ), .op(n11268) );
  nand2_1 U14173 ( .ip1(n11855), .ip2(\cache_data_B[2][48] ), .op(n11267) );
  nand2_1 U14174 ( .ip1(n12458), .ip2(\cache_data_B[6][48] ), .op(n11266) );
  nand2_1 U14175 ( .ip1(n10702), .ip2(\cache_data_B[7][48] ), .op(n11265) );
  nand4_1 U14176 ( .ip1(n11268), .ip2(n11267), .ip3(n11266), .ip4(n11265), 
        .op(n11269) );
  not_ab_or_c_or_d U14177 ( .ip1(\cache_data_B[0][48] ), .ip2(n12297), .ip3(
        n11270), .ip4(n11269), .op(n11272) );
  nand2_1 U14178 ( .ip1(n11296), .ip2(\cache_data_B[5][48] ), .op(n11271) );
  nand3_1 U14179 ( .ip1(n11273), .ip2(n11272), .ip3(n11271), .op(n12893) );
  nand2_1 U14180 ( .ip1(n12563), .ip2(n12893), .op(n11285) );
  nand2_1 U14181 ( .ip1(n11946), .ip2(\cache_data_A[1][112] ), .op(n11283) );
  and2_1 U14182 ( .ip1(n12194), .ip2(\cache_data_A[4][112] ), .op(n11279) );
  nand2_1 U14183 ( .ip1(n11855), .ip2(\cache_data_A[2][112] ), .op(n11277) );
  nand2_1 U14184 ( .ip1(n12410), .ip2(\cache_data_A[3][112] ), .op(n11276) );
  nand2_1 U14185 ( .ip1(n10702), .ip2(\cache_data_A[7][112] ), .op(n11275) );
  nand2_1 U14186 ( .ip1(n11780), .ip2(\cache_data_A[6][112] ), .op(n11274) );
  nand4_1 U14187 ( .ip1(n11277), .ip2(n11276), .ip3(n11275), .ip4(n11274), 
        .op(n11278) );
  not_ab_or_c_or_d U14188 ( .ip1(\cache_data_A[0][112] ), .ip2(n12357), .ip3(
        n11279), .ip4(n11278), .op(n11282) );
  nand2_1 U14189 ( .ip1(n11280), .ip2(\cache_data_A[5][112] ), .op(n11281) );
  nand3_1 U14190 ( .ip1(n11283), .ip2(n11282), .ip3(n11281), .op(n12895) );
  nand2_1 U14191 ( .ip1(n12509), .ip2(n12895), .op(n11284) );
  nand4_1 U14192 ( .ip1(n11287), .ip2(n11286), .ip3(n11285), .ip4(n11284), 
        .op(n11288) );
  not_ab_or_c_or_d U14193 ( .ip1(n12580), .ip2(n12890), .ip3(n11289), .ip4(
        n11288), .op(n11301) );
  nand2_1 U14194 ( .ip1(\cache_data_A[7][48] ), .ip2(n12552), .op(n11299) );
  and2_1 U14195 ( .ip1(n12476), .ip2(\cache_data_A[4][48] ), .op(n11295) );
  nand2_1 U14196 ( .ip1(n12321), .ip2(\cache_data_A[3][48] ), .op(n11293) );
  nand2_1 U14197 ( .ip1(n11911), .ip2(\cache_data_A[0][48] ), .op(n11292) );
  nand2_1 U14198 ( .ip1(n11946), .ip2(\cache_data_A[1][48] ), .op(n11291) );
  nand2_1 U14199 ( .ip1(n11780), .ip2(\cache_data_A[6][48] ), .op(n11290) );
  nand4_1 U14200 ( .ip1(n11293), .ip2(n11292), .ip3(n11291), .ip4(n11290), 
        .op(n11294) );
  not_ab_or_c_or_d U14201 ( .ip1(\cache_data_A[2][48] ), .ip2(n12546), .ip3(
        n11295), .ip4(n11294), .op(n11298) );
  nand2_1 U14202 ( .ip1(n11296), .ip2(\cache_data_A[5][48] ), .op(n11297) );
  nand3_1 U14203 ( .ip1(n11299), .ip2(n11298), .ip3(n11297), .op(n12894) );
  nand2_1 U14204 ( .ip1(n12595), .ip2(n12894), .op(n11300) );
  nand3_1 U14205 ( .ip1(n11302), .ip2(n11301), .ip3(n11300), .op(n11303) );
  mux2_1 U14206 ( .ip1(N4156), .ip2(n11303), .s(n11472), .op(n5304) );
  nand2_1 U14207 ( .ip1(n12552), .ip2(\cache_data_A[7][113] ), .op(n11314) );
  and2_1 U14208 ( .ip1(n12321), .ip2(\cache_data_A[3][113] ), .op(n11310) );
  nand2_1 U14209 ( .ip1(n12204), .ip2(\cache_data_A[0][113] ), .op(n11308) );
  nand2_1 U14210 ( .ip1(n11304), .ip2(\cache_data_A[5][113] ), .op(n11307) );
  nand2_1 U14211 ( .ip1(n11324), .ip2(\cache_data_A[4][113] ), .op(n11306) );
  nand2_1 U14212 ( .ip1(n11855), .ip2(\cache_data_A[2][113] ), .op(n11305) );
  nand4_1 U14213 ( .ip1(n11308), .ip2(n11307), .ip3(n11306), .ip4(n11305), 
        .op(n11309) );
  not_ab_or_c_or_d U14214 ( .ip1(\cache_data_A[6][113] ), .ip2(n12551), .ip3(
        n11310), .ip4(n11309), .op(n11313) );
  nand2_1 U14215 ( .ip1(n11311), .ip2(\cache_data_A[1][113] ), .op(n11312) );
  nand3_1 U14216 ( .ip1(n11314), .ip2(n11313), .ip3(n11312), .op(n12908) );
  nand2_1 U14217 ( .ip1(n12509), .ip2(n12908), .op(n11388) );
  nand2_1 U14218 ( .ip1(n12486), .ip2(\cache_data_A[2][17] ), .op(n11323) );
  and2_1 U14219 ( .ip1(n11946), .ip2(\cache_data_A[1][17] ), .op(n11320) );
  nand2_1 U14220 ( .ip1(n12591), .ip2(\cache_data_A[3][17] ), .op(n11318) );
  nand2_1 U14221 ( .ip1(n12584), .ip2(\cache_data_A[4][17] ), .op(n11317) );
  nand2_1 U14222 ( .ip1(n12458), .ip2(\cache_data_A[6][17] ), .op(n11316) );
  nand2_1 U14223 ( .ip1(n11911), .ip2(\cache_data_A[0][17] ), .op(n11315) );
  nand4_1 U14224 ( .ip1(n11318), .ip2(n11317), .ip3(n11316), .ip4(n11315), 
        .op(n11319) );
  not_ab_or_c_or_d U14225 ( .ip1(\cache_data_A[7][17] ), .ip2(n12278), .ip3(
        n11320), .ip4(n11319), .op(n11322) );
  nand2_1 U14226 ( .ip1(n12582), .ip2(\cache_data_A[5][17] ), .op(n11321) );
  nand3_1 U14227 ( .ip1(n11323), .ip2(n11322), .ip3(n11321), .op(n12911) );
  nand2_1 U14228 ( .ip1(n11780), .ip2(\cache_data_A[6][81] ), .op(n11328) );
  nand2_1 U14229 ( .ip1(n10575), .ip2(\cache_data_A[7][81] ), .op(n11327) );
  nand2_1 U14230 ( .ip1(n11946), .ip2(\cache_data_A[1][81] ), .op(n11326) );
  nand2_1 U14231 ( .ip1(n11324), .ip2(\cache_data_A[4][81] ), .op(n11325) );
  nand4_1 U14232 ( .ip1(n11328), .ip2(n11327), .ip3(n11326), .ip4(n11325), 
        .op(n11334) );
  nand2_1 U14233 ( .ip1(n12410), .ip2(\cache_data_A[3][81] ), .op(n11332) );
  nand2_1 U14234 ( .ip1(n12204), .ip2(\cache_data_A[0][81] ), .op(n11331) );
  nand2_1 U14235 ( .ip1(n11855), .ip2(\cache_data_A[2][81] ), .op(n11330) );
  nand2_1 U14236 ( .ip1(n12256), .ip2(\cache_data_A[5][81] ), .op(n11329) );
  nand4_1 U14237 ( .ip1(n11332), .ip2(n11331), .ip3(n11330), .ip4(n11329), 
        .op(n11333) );
  nor2_1 U14238 ( .ip1(n11334), .ip2(n11333), .op(n12909) );
  nor2_1 U14239 ( .ip1(n12909), .ip2(n12529), .op(n11376) );
  nand2_1 U14240 ( .ip1(n11780), .ip2(\cache_data_B[6][113] ), .op(n11343) );
  and2_1 U14241 ( .ip1(n11280), .ip2(\cache_data_B[5][113] ), .op(n11340) );
  nand2_1 U14242 ( .ip1(n12486), .ip2(\cache_data_B[2][113] ), .op(n11338) );
  nand2_1 U14243 ( .ip1(n12559), .ip2(\cache_data_B[3][113] ), .op(n11337) );
  nand2_1 U14244 ( .ip1(n12054), .ip2(\cache_data_B[4][113] ), .op(n11336) );
  nand2_1 U14245 ( .ip1(n12552), .ip2(\cache_data_B[7][113] ), .op(n11335) );
  nand4_1 U14246 ( .ip1(n11338), .ip2(n11337), .ip3(n11336), .ip4(n11335), 
        .op(n11339) );
  not_ab_or_c_or_d U14247 ( .ip1(n12297), .ip2(\cache_data_B[0][113] ), .ip3(
        n11340), .ip4(n11339), .op(n11342) );
  nand2_1 U14248 ( .ip1(n11946), .ip2(\cache_data_B[1][113] ), .op(n11341) );
  nand3_1 U14249 ( .ip1(n11343), .ip2(n11342), .ip3(n11341), .op(n12921) );
  nand2_1 U14250 ( .ip1(n12573), .ip2(n12921), .op(n11374) );
  nand2_1 U14251 ( .ip1(\cache_data_B[0][81] ), .ip2(n12204), .op(n11352) );
  and2_1 U14252 ( .ip1(n12371), .ip2(\cache_data_B[6][81] ), .op(n11349) );
  nand2_1 U14253 ( .ip1(n11946), .ip2(\cache_data_B[1][81] ), .op(n11347) );
  nand2_1 U14254 ( .ip1(n12591), .ip2(\cache_data_B[3][81] ), .op(n11346) );
  nand2_1 U14255 ( .ip1(n12054), .ip2(\cache_data_B[4][81] ), .op(n11345) );
  nand2_1 U14256 ( .ip1(n11855), .ip2(\cache_data_B[2][81] ), .op(n11344) );
  nand4_1 U14257 ( .ip1(n11347), .ip2(n11346), .ip3(n11345), .ip4(n11344), 
        .op(n11348) );
  not_ab_or_c_or_d U14258 ( .ip1(n12278), .ip2(\cache_data_B[7][81] ), .ip3(
        n11349), .ip4(n11348), .op(n11351) );
  nand2_1 U14259 ( .ip1(n11280), .ip2(\cache_data_B[5][81] ), .op(n11350) );
  nand3_1 U14260 ( .ip1(n11352), .ip2(n11351), .ip3(n11350), .op(n12912) );
  nand2_1 U14261 ( .ip1(n12580), .ip2(n12912), .op(n11373) );
  nand2_1 U14262 ( .ip1(\cache_data_B[6][17] ), .ip2(n12371), .op(n11361) );
  and2_1 U14263 ( .ip1(n12476), .ip2(\cache_data_B[4][17] ), .op(n11358) );
  nand2_1 U14264 ( .ip1(n12486), .ip2(\cache_data_B[2][17] ), .op(n11356) );
  buf_1 U14265 ( .ip(n11724), .op(n12242) );
  nand2_1 U14266 ( .ip1(n12242), .ip2(\cache_data_B[1][17] ), .op(n11355) );
  nand2_1 U14267 ( .ip1(n12204), .ip2(\cache_data_B[0][17] ), .op(n11354) );
  nand2_1 U14268 ( .ip1(n11236), .ip2(\cache_data_B[5][17] ), .op(n11353) );
  nand4_1 U14269 ( .ip1(n11356), .ip2(n11355), .ip3(n11354), .ip4(n11353), 
        .op(n11357) );
  not_ab_or_c_or_d U14270 ( .ip1(\cache_data_B[7][17] ), .ip2(n12278), .ip3(
        n11358), .ip4(n11357), .op(n11360) );
  nand2_1 U14271 ( .ip1(n12321), .ip2(\cache_data_B[3][17] ), .op(n11359) );
  nand3_1 U14272 ( .ip1(n11361), .ip2(n11360), .ip3(n11359), .op(n12913) );
  nand2_1 U14273 ( .ip1(n12539), .ip2(n12913), .op(n11372) );
  nand2_1 U14274 ( .ip1(\cache_data_A[3][49] ), .ip2(n12410), .op(n11370) );
  and2_1 U14275 ( .ip1(n10686), .ip2(\cache_data_A[1][49] ), .op(n11367) );
  nand2_1 U14276 ( .ip1(n12551), .ip2(\cache_data_A[6][49] ), .op(n11365) );
  nand2_1 U14277 ( .ip1(n12584), .ip2(\cache_data_A[4][49] ), .op(n11364) );
  nand2_1 U14278 ( .ip1(n12486), .ip2(\cache_data_A[2][49] ), .op(n11363) );
  nand2_1 U14279 ( .ip1(n11911), .ip2(\cache_data_A[0][49] ), .op(n11362) );
  nand4_1 U14280 ( .ip1(n11365), .ip2(n11364), .ip3(n11363), .ip4(n11362), 
        .op(n11366) );
  not_ab_or_c_or_d U14281 ( .ip1(n12278), .ip2(\cache_data_A[7][49] ), .ip3(
        n11367), .ip4(n11366), .op(n11369) );
  nand2_1 U14282 ( .ip1(n11280), .ip2(\cache_data_A[5][49] ), .op(n11368) );
  nand3_1 U14283 ( .ip1(n11370), .ip2(n11369), .ip3(n11368), .op(n12910) );
  nand2_1 U14284 ( .ip1(n12595), .ip2(n12910), .op(n11371) );
  nand4_1 U14285 ( .ip1(n11374), .ip2(n11373), .ip3(n11372), .ip4(n11371), 
        .op(n11375) );
  not_ab_or_c_or_d U14286 ( .ip1(n12550), .ip2(n12911), .ip3(n11376), .ip4(
        n11375), .op(n11387) );
  nand2_1 U14287 ( .ip1(n12204), .ip2(\cache_data_B[0][49] ), .op(n11385) );
  and2_1 U14288 ( .ip1(n12458), .ip2(\cache_data_B[6][49] ), .op(n11382) );
  nand2_1 U14289 ( .ip1(n8060), .ip2(\cache_data_B[3][49] ), .op(n11380) );
  nand2_1 U14290 ( .ip1(n10575), .ip2(\cache_data_B[7][49] ), .op(n11379) );
  nand2_1 U14291 ( .ip1(n11724), .ip2(\cache_data_B[1][49] ), .op(n11378) );
  nand2_1 U14292 ( .ip1(n11156), .ip2(\cache_data_B[4][49] ), .op(n11377) );
  nand4_1 U14293 ( .ip1(n11380), .ip2(n11379), .ip3(n11378), .ip4(n11377), 
        .op(n11381) );
  not_ab_or_c_or_d U14294 ( .ip1(n12546), .ip2(\cache_data_B[2][49] ), .ip3(
        n11382), .ip4(n11381), .op(n11384) );
  nand2_1 U14295 ( .ip1(n12118), .ip2(\cache_data_B[5][49] ), .op(n11383) );
  nand3_1 U14296 ( .ip1(n11385), .ip2(n11384), .ip3(n11383), .op(n12920) );
  nand2_1 U14297 ( .ip1(n12563), .ip2(n12920), .op(n11386) );
  nand3_1 U14298 ( .ip1(n11388), .ip2(n11387), .ip3(n11386), .op(n11389) );
  mux2_1 U14299 ( .ip1(N4153), .ip2(n11389), .s(n11472), .op(n5303) );
  nand2_1 U14300 ( .ip1(n11911), .ip2(\cache_data_B[0][50] ), .op(n11398) );
  and2_1 U14301 ( .ip1(n11296), .ip2(\cache_data_B[5][50] ), .op(n11395) );
  nand2_1 U14302 ( .ip1(n11780), .ip2(\cache_data_B[6][50] ), .op(n11393) );
  nand2_1 U14303 ( .ip1(n11057), .ip2(\cache_data_B[7][50] ), .op(n11392) );
  nand2_1 U14304 ( .ip1(n11855), .ip2(\cache_data_B[2][50] ), .op(n11391) );
  nand2_1 U14305 ( .ip1(n8060), .ip2(\cache_data_B[3][50] ), .op(n11390) );
  nand4_1 U14306 ( .ip1(n11393), .ip2(n11392), .ip3(n11391), .ip4(n11390), 
        .op(n11394) );
  not_ab_or_c_or_d U14307 ( .ip1(n11946), .ip2(\cache_data_B[1][50] ), .ip3(
        n11395), .ip4(n11394), .op(n11397) );
  nand2_1 U14308 ( .ip1(n12584), .ip2(\cache_data_B[4][50] ), .op(n11396) );
  nand3_1 U14309 ( .ip1(n11398), .ip2(n11397), .ip3(n11396), .op(n12929) );
  nand2_1 U14310 ( .ip1(n12563), .ip2(n12929), .op(n11471) );
  nand2_1 U14311 ( .ip1(\cache_data_B[7][82] ), .ip2(n12552), .op(n11407) );
  and2_1 U14312 ( .ip1(n11304), .ip2(\cache_data_B[5][82] ), .op(n11404) );
  nand2_1 U14313 ( .ip1(n12204), .ip2(\cache_data_B[0][82] ), .op(n11402) );
  nand2_1 U14314 ( .ip1(n11780), .ip2(\cache_data_B[6][82] ), .op(n11401) );
  nand2_1 U14315 ( .ip1(n12486), .ip2(\cache_data_B[2][82] ), .op(n11400) );
  nand2_1 U14316 ( .ip1(n12242), .ip2(\cache_data_B[1][82] ), .op(n11399) );
  nand4_1 U14317 ( .ip1(n11402), .ip2(n11401), .ip3(n11400), .ip4(n11399), 
        .op(n11403) );
  not_ab_or_c_or_d U14318 ( .ip1(\cache_data_B[4][82] ), .ip2(n12476), .ip3(
        n11404), .ip4(n11403), .op(n11406) );
  nand2_1 U14319 ( .ip1(n12321), .ip2(\cache_data_B[3][82] ), .op(n11405) );
  nand3_1 U14320 ( .ip1(n11407), .ip2(n11406), .ip3(n11405), .op(n12928) );
  nand2_1 U14321 ( .ip1(n12321), .ip2(\cache_data_A[3][82] ), .op(n11411) );
  nand2_1 U14322 ( .ip1(n12371), .ip2(\cache_data_A[6][82] ), .op(n11410) );
  nand2_1 U14323 ( .ip1(n12204), .ip2(\cache_data_A[0][82] ), .op(n11409) );
  nand2_1 U14324 ( .ip1(n12194), .ip2(\cache_data_A[4][82] ), .op(n11408) );
  nand4_1 U14325 ( .ip1(n11411), .ip2(n11410), .ip3(n11409), .ip4(n11408), 
        .op(n11417) );
  nand2_1 U14326 ( .ip1(n12118), .ip2(\cache_data_A[5][82] ), .op(n11415) );
  nand2_1 U14327 ( .ip1(n10575), .ip2(\cache_data_A[7][82] ), .op(n11414) );
  nand2_1 U14328 ( .ip1(n11855), .ip2(\cache_data_A[2][82] ), .op(n11413) );
  nand2_1 U14329 ( .ip1(n12147), .ip2(\cache_data_A[1][82] ), .op(n11412) );
  nand4_1 U14330 ( .ip1(n11415), .ip2(n11414), .ip3(n11413), .ip4(n11412), 
        .op(n11416) );
  nor2_1 U14331 ( .ip1(n11417), .ip2(n11416), .op(n12927) );
  nor2_1 U14332 ( .ip1(n12927), .ip2(n12529), .op(n11459) );
  nand2_1 U14333 ( .ip1(\cache_data_B[4][114] ), .ip2(n12194), .op(n11426) );
  and2_1 U14334 ( .ip1(n12321), .ip2(\cache_data_B[3][114] ), .op(n11423) );
  nand2_1 U14335 ( .ip1(n11911), .ip2(\cache_data_B[0][114] ), .op(n11421) );
  nand2_1 U14336 ( .ip1(n12486), .ip2(\cache_data_B[2][114] ), .op(n11420) );
  nand2_1 U14337 ( .ip1(n11236), .ip2(\cache_data_B[5][114] ), .op(n11419) );
  nand2_1 U14338 ( .ip1(n12468), .ip2(\cache_data_B[7][114] ), .op(n11418) );
  nand4_1 U14339 ( .ip1(n11421), .ip2(n11420), .ip3(n11419), .ip4(n11418), 
        .op(n11422) );
  not_ab_or_c_or_d U14340 ( .ip1(n12551), .ip2(\cache_data_B[6][114] ), .ip3(
        n11423), .ip4(n11422), .op(n11425) );
  nand2_1 U14341 ( .ip1(n11724), .ip2(\cache_data_B[1][114] ), .op(n11424) );
  nand3_1 U14342 ( .ip1(n11426), .ip2(n11425), .ip3(n11424), .op(n12939) );
  nand2_1 U14343 ( .ip1(n12573), .ip2(n12939), .op(n11457) );
  nand2_1 U14344 ( .ip1(n11855), .ip2(\cache_data_A[2][114] ), .op(n11435) );
  and2_1 U14345 ( .ip1(n11946), .ip2(\cache_data_A[1][114] ), .op(n11432) );
  nand2_1 U14346 ( .ip1(n12591), .ip2(\cache_data_A[3][114] ), .op(n11430) );
  nand2_1 U14347 ( .ip1(n12194), .ip2(\cache_data_A[4][114] ), .op(n11429) );
  nand2_1 U14348 ( .ip1(n12204), .ip2(\cache_data_A[0][114] ), .op(n11428) );
  nand2_1 U14349 ( .ip1(n12118), .ip2(\cache_data_A[5][114] ), .op(n11427) );
  nand4_1 U14350 ( .ip1(n11430), .ip2(n11429), .ip3(n11428), .ip4(n11427), 
        .op(n11431) );
  not_ab_or_c_or_d U14351 ( .ip1(\cache_data_A[7][114] ), .ip2(n12278), .ip3(
        n11432), .ip4(n11431), .op(n11434) );
  nand2_1 U14352 ( .ip1(n11780), .ip2(\cache_data_A[6][114] ), .op(n11433) );
  nand3_1 U14353 ( .ip1(n11435), .ip2(n11434), .ip3(n11433), .op(n12930) );
  nand2_1 U14354 ( .ip1(n12509), .ip2(n12930), .op(n11456) );
  nand2_1 U14355 ( .ip1(n12204), .ip2(\cache_data_A[0][18] ), .op(n11444) );
  and2_1 U14356 ( .ip1(n12256), .ip2(\cache_data_A[5][18] ), .op(n11441) );
  nand2_1 U14357 ( .ip1(n12486), .ip2(\cache_data_A[2][18] ), .op(n11439) );
  nand2_1 U14358 ( .ip1(n12429), .ip2(\cache_data_A[6][18] ), .op(n11438) );
  nand2_1 U14359 ( .ip1(n12147), .ip2(\cache_data_A[1][18] ), .op(n11437) );
  nand2_1 U14360 ( .ip1(n11324), .ip2(\cache_data_A[4][18] ), .op(n11436) );
  nand4_1 U14361 ( .ip1(n11439), .ip2(n11438), .ip3(n11437), .ip4(n11436), 
        .op(n11440) );
  not_ab_or_c_or_d U14362 ( .ip1(\cache_data_A[3][18] ), .ip2(n12559), .ip3(
        n11441), .ip4(n11440), .op(n11443) );
  nand2_1 U14363 ( .ip1(n11057), .ip2(\cache_data_A[7][18] ), .op(n11442) );
  nand3_1 U14364 ( .ip1(n11444), .ip2(n11443), .ip3(n11442), .op(n12938) );
  nand2_1 U14365 ( .ip1(n12550), .ip2(n12938), .op(n11455) );
  nand2_1 U14366 ( .ip1(n12410), .ip2(\cache_data_A[3][50] ), .op(n11453) );
  and2_1 U14367 ( .ip1(n11946), .ip2(\cache_data_A[1][50] ), .op(n11450) );
  nand2_1 U14368 ( .ip1(n11855), .ip2(\cache_data_A[2][50] ), .op(n11448) );
  nand2_1 U14369 ( .ip1(n12584), .ip2(\cache_data_A[4][50] ), .op(n11447) );
  nand2_1 U14370 ( .ip1(n11057), .ip2(\cache_data_A[7][50] ), .op(n11446) );
  nand2_1 U14371 ( .ip1(n11780), .ip2(\cache_data_A[6][50] ), .op(n11445) );
  nand4_1 U14372 ( .ip1(n11448), .ip2(n11447), .ip3(n11446), .ip4(n11445), 
        .op(n11449) );
  not_ab_or_c_or_d U14373 ( .ip1(\cache_data_A[0][50] ), .ip2(n12297), .ip3(
        n11450), .ip4(n11449), .op(n11452) );
  nand2_1 U14374 ( .ip1(n12256), .ip2(\cache_data_A[5][50] ), .op(n11451) );
  nand3_1 U14375 ( .ip1(n11453), .ip2(n11452), .ip3(n11451), .op(n12931) );
  nand2_1 U14376 ( .ip1(n12595), .ip2(n12931), .op(n11454) );
  nand4_1 U14377 ( .ip1(n11457), .ip2(n11456), .ip3(n11455), .ip4(n11454), 
        .op(n11458) );
  not_ab_or_c_or_d U14378 ( .ip1(n12580), .ip2(n12928), .ip3(n11459), .ip4(
        n11458), .op(n11470) );
  nand2_1 U14379 ( .ip1(n11911), .ip2(\cache_data_B[0][18] ), .op(n11468) );
  and2_1 U14380 ( .ip1(n12147), .ip2(\cache_data_B[1][18] ), .op(n11465) );
  nand2_1 U14381 ( .ip1(n12584), .ip2(\cache_data_B[4][18] ), .op(n11463) );
  nand2_1 U14382 ( .ip1(n12410), .ip2(\cache_data_B[3][18] ), .op(n11462) );
  nand2_1 U14383 ( .ip1(n10575), .ip2(\cache_data_B[7][18] ), .op(n11461) );
  nand2_1 U14384 ( .ip1(n12256), .ip2(\cache_data_B[5][18] ), .op(n11460) );
  nand4_1 U14385 ( .ip1(n11463), .ip2(n11462), .ip3(n11461), .ip4(n11460), 
        .op(n11464) );
  not_ab_or_c_or_d U14386 ( .ip1(\cache_data_B[2][18] ), .ip2(n12475), .ip3(
        n11465), .ip4(n11464), .op(n11467) );
  nand2_1 U14387 ( .ip1(n11780), .ip2(\cache_data_B[6][18] ), .op(n11466) );
  nand3_1 U14388 ( .ip1(n11468), .ip2(n11467), .ip3(n11466), .op(n12926) );
  nand2_1 U14389 ( .ip1(n12539), .ip2(n12926), .op(n11469) );
  nand3_1 U14390 ( .ip1(n11471), .ip2(n11470), .ip3(n11469), .op(n11473) );
  mux2_1 U14391 ( .ip1(N4150), .ip2(n11473), .s(n11472), .op(n5302) );
  nand2_1 U14392 ( .ip1(\cache_data_A[3][51] ), .ip2(n12410), .op(n11482) );
  and2_1 U14393 ( .ip1(n12118), .ip2(\cache_data_A[5][51] ), .op(n11479) );
  nand2_1 U14394 ( .ip1(n11780), .ip2(\cache_data_A[6][51] ), .op(n11477) );
  nand2_1 U14395 ( .ip1(n11911), .ip2(\cache_data_A[0][51] ), .op(n11476) );
  nand2_1 U14396 ( .ip1(n12468), .ip2(\cache_data_A[7][51] ), .op(n11475) );
  nand2_1 U14397 ( .ip1(n11855), .ip2(\cache_data_A[2][51] ), .op(n11474) );
  nand4_1 U14398 ( .ip1(n11477), .ip2(n11476), .ip3(n11475), .ip4(n11474), 
        .op(n11478) );
  not_ab_or_c_or_d U14399 ( .ip1(n11156), .ip2(\cache_data_A[4][51] ), .ip3(
        n11479), .ip4(n11478), .op(n11481) );
  nand2_1 U14400 ( .ip1(n11724), .ip2(\cache_data_A[1][51] ), .op(n11480) );
  nand3_1 U14401 ( .ip1(n11482), .ip2(n11481), .ip3(n11480), .op(n12957) );
  nand2_1 U14402 ( .ip1(n12595), .ip2(n12957), .op(n11556) );
  nand2_1 U14403 ( .ip1(\cache_data_A[0][19] ), .ip2(n12204), .op(n11491) );
  and2_1 U14404 ( .ip1(n12582), .ip2(\cache_data_A[5][19] ), .op(n11488) );
  nand2_1 U14405 ( .ip1(n12147), .ip2(\cache_data_A[1][19] ), .op(n11486) );
  nand2_1 U14406 ( .ip1(n12591), .ip2(\cache_data_A[3][19] ), .op(n11485) );
  nand2_1 U14407 ( .ip1(n12429), .ip2(\cache_data_A[6][19] ), .op(n11484) );
  nand2_1 U14408 ( .ip1(n11855), .ip2(\cache_data_A[2][19] ), .op(n11483) );
  nand4_1 U14409 ( .ip1(n11486), .ip2(n11485), .ip3(n11484), .ip4(n11483), 
        .op(n11487) );
  not_ab_or_c_or_d U14410 ( .ip1(\cache_data_A[7][19] ), .ip2(n10702), .ip3(
        n11488), .ip4(n11487), .op(n11490) );
  nand2_1 U14411 ( .ip1(n12584), .ip2(\cache_data_A[4][19] ), .op(n11489) );
  nand3_1 U14412 ( .ip1(n11491), .ip2(n11490), .ip3(n11489), .op(n12949) );
  nand2_1 U14413 ( .ip1(n11911), .ip2(\cache_data_A[0][83] ), .op(n11495) );
  nand2_1 U14414 ( .ip1(n11780), .ip2(\cache_data_A[6][83] ), .op(n11494) );
  nand2_1 U14415 ( .ip1(n12552), .ip2(\cache_data_A[7][83] ), .op(n11493) );
  nand2_1 U14416 ( .ip1(n12476), .ip2(\cache_data_A[4][83] ), .op(n11492) );
  nand4_1 U14417 ( .ip1(n11495), .ip2(n11494), .ip3(n11493), .ip4(n11492), 
        .op(n11501) );
  nand2_1 U14418 ( .ip1(n11855), .ip2(\cache_data_A[2][83] ), .op(n11499) );
  nand2_1 U14419 ( .ip1(n12410), .ip2(\cache_data_A[3][83] ), .op(n11498) );
  nand2_1 U14420 ( .ip1(n11724), .ip2(\cache_data_A[1][83] ), .op(n11497) );
  nand2_1 U14421 ( .ip1(n11280), .ip2(\cache_data_A[5][83] ), .op(n11496) );
  nand4_1 U14422 ( .ip1(n11499), .ip2(n11498), .ip3(n11497), .ip4(n11496), 
        .op(n11500) );
  nor2_1 U14423 ( .ip1(n11501), .ip2(n11500), .op(n12945) );
  nor2_1 U14424 ( .ip1(n12945), .ip2(n12529), .op(n11544) );
  nand2_1 U14425 ( .ip1(n12410), .ip2(\cache_data_A[3][115] ), .op(n11510) );
  and2_1 U14426 ( .ip1(n10686), .ip2(\cache_data_A[1][115] ), .op(n11507) );
  nand2_1 U14427 ( .ip1(n11780), .ip2(\cache_data_A[6][115] ), .op(n11505) );
  nand2_1 U14428 ( .ip1(n11855), .ip2(\cache_data_A[2][115] ), .op(n11504) );
  nand2_1 U14429 ( .ip1(n11911), .ip2(\cache_data_A[0][115] ), .op(n11503) );
  nand2_1 U14430 ( .ip1(n12118), .ip2(\cache_data_A[5][115] ), .op(n11502) );
  nand4_1 U14431 ( .ip1(n11505), .ip2(n11504), .ip3(n11503), .ip4(n11502), 
        .op(n11506) );
  not_ab_or_c_or_d U14432 ( .ip1(\cache_data_A[7][115] ), .ip2(n12278), .ip3(
        n11507), .ip4(n11506), .op(n11509) );
  nand2_1 U14433 ( .ip1(n12584), .ip2(\cache_data_A[4][115] ), .op(n11508) );
  nand3_1 U14434 ( .ip1(n11510), .ip2(n11509), .ip3(n11508), .op(n12947) );
  nand2_1 U14435 ( .ip1(n12509), .ip2(n12947), .op(n11542) );
  nand2_1 U14436 ( .ip1(n11911), .ip2(\cache_data_B[0][83] ), .op(n11519) );
  and2_1 U14437 ( .ip1(n12476), .ip2(\cache_data_B[4][83] ), .op(n11516) );
  nand2_1 U14438 ( .ip1(n11855), .ip2(\cache_data_B[2][83] ), .op(n11514) );
  nand2_1 U14439 ( .ip1(n12147), .ip2(\cache_data_B[1][83] ), .op(n11513) );
  nand2_1 U14440 ( .ip1(n12118), .ip2(\cache_data_B[5][83] ), .op(n11512) );
  nand2_1 U14441 ( .ip1(n12581), .ip2(\cache_data_B[7][83] ), .op(n11511) );
  nand4_1 U14442 ( .ip1(n11514), .ip2(n11513), .ip3(n11512), .ip4(n11511), 
        .op(n11515) );
  not_ab_or_c_or_d U14443 ( .ip1(\cache_data_B[6][83] ), .ip2(n12551), .ip3(
        n11516), .ip4(n11515), .op(n11518) );
  nand2_1 U14444 ( .ip1(n8060), .ip2(\cache_data_B[3][83] ), .op(n11517) );
  nand3_1 U14445 ( .ip1(n11519), .ip2(n11518), .ip3(n11517), .op(n12944) );
  nand2_1 U14446 ( .ip1(n12580), .ip2(n12944), .op(n11541) );
  nand2_1 U14447 ( .ip1(n11911), .ip2(\cache_data_B[0][51] ), .op(n11528) );
  and2_1 U14448 ( .ip1(n12591), .ip2(\cache_data_B[3][51] ), .op(n11525) );
  nand2_1 U14449 ( .ip1(n12147), .ip2(\cache_data_B[1][51] ), .op(n11523) );
  nand2_1 U14450 ( .ip1(n11236), .ip2(\cache_data_B[5][51] ), .op(n11522) );
  nand2_1 U14451 ( .ip1(n11855), .ip2(\cache_data_B[2][51] ), .op(n11521) );
  nand2_1 U14452 ( .ip1(n12584), .ip2(\cache_data_B[4][51] ), .op(n11520) );
  nand4_1 U14453 ( .ip1(n11523), .ip2(n11522), .ip3(n11521), .ip4(n11520), 
        .op(n11524) );
  not_ab_or_c_or_d U14454 ( .ip1(n12278), .ip2(\cache_data_B[7][51] ), .ip3(
        n11525), .ip4(n11524), .op(n11527) );
  nand2_1 U14455 ( .ip1(n11780), .ip2(\cache_data_B[6][51] ), .op(n11526) );
  nand3_1 U14456 ( .ip1(n11528), .ip2(n11527), .ip3(n11526), .op(n12948) );
  nand2_1 U14457 ( .ip1(n12563), .ip2(n12948), .op(n11540) );
  nand2_1 U14458 ( .ip1(\cache_data_B[2][115] ), .ip2(n12486), .op(n11538) );
  and2_1 U14459 ( .ip1(n12476), .ip2(\cache_data_B[4][115] ), .op(n11534) );
  nand2_1 U14460 ( .ip1(n11780), .ip2(\cache_data_B[6][115] ), .op(n11532) );
  nand2_1 U14461 ( .ip1(n11911), .ip2(\cache_data_B[0][115] ), .op(n11531) );
  nand2_1 U14462 ( .ip1(n10702), .ip2(\cache_data_B[7][115] ), .op(n11530) );
  nand2_1 U14463 ( .ip1(n12147), .ip2(\cache_data_B[1][115] ), .op(n11529) );
  nand4_1 U14464 ( .ip1(n11532), .ip2(n11531), .ip3(n11530), .ip4(n11529), 
        .op(n11533) );
  not_ab_or_c_or_d U14465 ( .ip1(\cache_data_B[3][115] ), .ip2(n11535), .ip3(
        n11534), .ip4(n11533), .op(n11537) );
  nand2_1 U14466 ( .ip1(n12256), .ip2(\cache_data_B[5][115] ), .op(n11536) );
  nand3_1 U14467 ( .ip1(n11538), .ip2(n11537), .ip3(n11536), .op(n12956) );
  nand2_1 U14468 ( .ip1(n12573), .ip2(n12956), .op(n11539) );
  nand4_1 U14469 ( .ip1(n11542), .ip2(n11541), .ip3(n11540), .ip4(n11539), 
        .op(n11543) );
  not_ab_or_c_or_d U14470 ( .ip1(n12550), .ip2(n12949), .ip3(n11544), .ip4(
        n11543), .op(n11555) );
  nand2_1 U14471 ( .ip1(n11724), .ip2(\cache_data_B[1][19] ), .op(n11553) );
  and2_1 U14472 ( .ip1(n12371), .ip2(\cache_data_B[6][19] ), .op(n11550) );
  nand2_1 U14473 ( .ip1(n12591), .ip2(\cache_data_B[3][19] ), .op(n11548) );
  nand2_1 U14474 ( .ip1(n11156), .ip2(\cache_data_B[4][19] ), .op(n11547) );
  nand2_1 U14475 ( .ip1(n11911), .ip2(\cache_data_B[0][19] ), .op(n11546) );
  nand2_1 U14476 ( .ip1(n11855), .ip2(\cache_data_B[2][19] ), .op(n11545) );
  nand4_1 U14477 ( .ip1(n11548), .ip2(n11547), .ip3(n11546), .ip4(n11545), 
        .op(n11549) );
  not_ab_or_c_or_d U14478 ( .ip1(\cache_data_B[7][19] ), .ip2(n12278), .ip3(
        n11550), .ip4(n11549), .op(n11552) );
  nand2_1 U14479 ( .ip1(n12256), .ip2(\cache_data_B[5][19] ), .op(n11551) );
  nand3_1 U14480 ( .ip1(n11553), .ip2(n11552), .ip3(n11551), .op(n12946) );
  nand2_1 U14481 ( .ip1(n12539), .ip2(n12946), .op(n11554) );
  nand3_1 U14482 ( .ip1(n11556), .ip2(n11555), .ip3(n11554), .op(n11557) );
  mux2_1 U14483 ( .ip1(N4147), .ip2(n11557), .s(n12599), .op(n5301) );
  nand2_1 U14484 ( .ip1(n12584), .ip2(\cache_data_A[4][20] ), .op(n11566) );
  and2_1 U14485 ( .ip1(n11296), .ip2(\cache_data_A[5][20] ), .op(n11563) );
  nand2_1 U14486 ( .ip1(n12581), .ip2(\cache_data_A[7][20] ), .op(n11561) );
  nand2_1 U14487 ( .ip1(n11855), .ip2(\cache_data_A[2][20] ), .op(n11560) );
  nand2_1 U14488 ( .ip1(n12410), .ip2(\cache_data_A[3][20] ), .op(n11559) );
  nand2_1 U14489 ( .ip1(n11780), .ip2(\cache_data_A[6][20] ), .op(n11558) );
  nand4_1 U14490 ( .ip1(n11561), .ip2(n11560), .ip3(n11559), .ip4(n11558), 
        .op(n11562) );
  not_ab_or_c_or_d U14491 ( .ip1(\cache_data_A[0][20] ), .ip2(n12297), .ip3(
        n11563), .ip4(n11562), .op(n11565) );
  nand2_1 U14492 ( .ip1(n11724), .ip2(\cache_data_A[1][20] ), .op(n11564) );
  nand3_1 U14493 ( .ip1(n11566), .ip2(n11565), .ip3(n11564), .op(n12962) );
  nand2_1 U14494 ( .ip1(n12550), .ip2(n12962), .op(n11639) );
  nand2_1 U14495 ( .ip1(\cache_data_B[2][52] ), .ip2(n12486), .op(n11575) );
  and2_1 U14496 ( .ip1(n12582), .ip2(\cache_data_B[5][52] ), .op(n11572) );
  nand2_1 U14497 ( .ip1(n10575), .ip2(\cache_data_B[7][52] ), .op(n11570) );
  nand2_1 U14498 ( .ip1(n8060), .ip2(\cache_data_B[3][52] ), .op(n11569) );
  nand2_1 U14499 ( .ip1(n12147), .ip2(\cache_data_B[1][52] ), .op(n11568) );
  nand2_1 U14500 ( .ip1(n11911), .ip2(\cache_data_B[0][52] ), .op(n11567) );
  nand4_1 U14501 ( .ip1(n11570), .ip2(n11569), .ip3(n11568), .ip4(n11567), 
        .op(n11571) );
  not_ab_or_c_or_d U14502 ( .ip1(n12551), .ip2(\cache_data_B[6][52] ), .ip3(
        n11572), .ip4(n11571), .op(n11574) );
  nand2_1 U14503 ( .ip1(n12476), .ip2(\cache_data_B[4][52] ), .op(n11573) );
  nand3_1 U14504 ( .ip1(n11575), .ip2(n11574), .ip3(n11573), .op(n12964) );
  nand2_1 U14505 ( .ip1(n12118), .ip2(\cache_data_A[5][84] ), .op(n11579) );
  nand2_1 U14506 ( .ip1(n11855), .ip2(\cache_data_A[2][84] ), .op(n11578) );
  nand2_1 U14507 ( .ip1(n10575), .ip2(\cache_data_A[7][84] ), .op(n11577) );
  nand2_1 U14508 ( .ip1(n11780), .ip2(\cache_data_A[6][84] ), .op(n11576) );
  nand4_1 U14509 ( .ip1(n11579), .ip2(n11578), .ip3(n11577), .ip4(n11576), 
        .op(n11585) );
  nand2_1 U14510 ( .ip1(n11911), .ip2(\cache_data_A[0][84] ), .op(n11583) );
  nand2_1 U14511 ( .ip1(n12584), .ip2(\cache_data_A[4][84] ), .op(n11582) );
  nand2_1 U14512 ( .ip1(n12410), .ip2(\cache_data_A[3][84] ), .op(n11581) );
  nand2_1 U14513 ( .ip1(n11724), .ip2(\cache_data_A[1][84] ), .op(n11580) );
  nand4_1 U14514 ( .ip1(n11583), .ip2(n11582), .ip3(n11581), .ip4(n11580), 
        .op(n11584) );
  nor2_1 U14515 ( .ip1(n11585), .ip2(n11584), .op(n12963) );
  nor2_1 U14516 ( .ip1(n12963), .ip2(n12529), .op(n11627) );
  nand2_1 U14517 ( .ip1(n11780), .ip2(\cache_data_B[6][84] ), .op(n11594) );
  and2_1 U14518 ( .ip1(n12591), .ip2(\cache_data_B[3][84] ), .op(n11591) );
  nand2_1 U14519 ( .ip1(n12242), .ip2(\cache_data_B[1][84] ), .op(n11589) );
  nand2_1 U14520 ( .ip1(n12054), .ip2(\cache_data_B[4][84] ), .op(n11588) );
  nand2_1 U14521 ( .ip1(n12581), .ip2(\cache_data_B[7][84] ), .op(n11587) );
  nand2_1 U14522 ( .ip1(n11911), .ip2(\cache_data_B[0][84] ), .op(n11586) );
  nand4_1 U14523 ( .ip1(n11589), .ip2(n11588), .ip3(n11587), .ip4(n11586), 
        .op(n11590) );
  not_ab_or_c_or_d U14524 ( .ip1(\cache_data_B[2][84] ), .ip2(n12546), .ip3(
        n11591), .ip4(n11590), .op(n11593) );
  nand2_1 U14525 ( .ip1(n12256), .ip2(\cache_data_B[5][84] ), .op(n11592) );
  nand3_1 U14526 ( .ip1(n11594), .ip2(n11593), .ip3(n11592), .op(n12975) );
  nand2_1 U14527 ( .ip1(n12580), .ip2(n12975), .op(n11625) );
  nand2_1 U14528 ( .ip1(\cache_data_B[7][116] ), .ip2(n12552), .op(n11603) );
  and2_1 U14529 ( .ip1(n12256), .ip2(\cache_data_B[5][116] ), .op(n11600) );
  nand2_1 U14530 ( .ip1(n11911), .ip2(\cache_data_B[0][116] ), .op(n11598) );
  nand2_1 U14531 ( .ip1(n12584), .ip2(\cache_data_B[4][116] ), .op(n11597) );
  nand2_1 U14532 ( .ip1(n12147), .ip2(\cache_data_B[1][116] ), .op(n11596) );
  nand2_1 U14533 ( .ip1(n11780), .ip2(\cache_data_B[6][116] ), .op(n11595) );
  nand4_1 U14534 ( .ip1(n11598), .ip2(n11597), .ip3(n11596), .ip4(n11595), 
        .op(n11599) );
  not_ab_or_c_or_d U14535 ( .ip1(n12546), .ip2(\cache_data_B[2][116] ), .ip3(
        n11600), .ip4(n11599), .op(n11602) );
  nand2_1 U14536 ( .ip1(n12410), .ip2(\cache_data_B[3][116] ), .op(n11601) );
  nand3_1 U14537 ( .ip1(n11603), .ip2(n11602), .ip3(n11601), .op(n12974) );
  nand2_1 U14538 ( .ip1(n12573), .ip2(n12974), .op(n11624) );
  nand2_1 U14539 ( .ip1(n11780), .ip2(\cache_data_A[6][116] ), .op(n11612) );
  and2_1 U14540 ( .ip1(n11946), .ip2(\cache_data_A[1][116] ), .op(n11609) );
  nand2_1 U14541 ( .ip1(n11911), .ip2(\cache_data_A[0][116] ), .op(n11607) );
  nand2_1 U14542 ( .ip1(n12584), .ip2(\cache_data_A[4][116] ), .op(n11606) );
  nand2_1 U14543 ( .ip1(n12410), .ip2(\cache_data_A[3][116] ), .op(n11605) );
  nand2_1 U14544 ( .ip1(n11855), .ip2(\cache_data_A[2][116] ), .op(n11604) );
  nand4_1 U14545 ( .ip1(n11607), .ip2(n11606), .ip3(n11605), .ip4(n11604), 
        .op(n11608) );
  not_ab_or_c_or_d U14546 ( .ip1(\cache_data_A[7][116] ), .ip2(n12278), .ip3(
        n11609), .ip4(n11608), .op(n11611) );
  nand2_1 U14547 ( .ip1(n12118), .ip2(\cache_data_A[5][116] ), .op(n11610) );
  nand3_1 U14548 ( .ip1(n11612), .ip2(n11611), .ip3(n11610), .op(n12966) );
  nand2_1 U14549 ( .ip1(n12509), .ip2(n12966), .op(n11623) );
  nand2_1 U14550 ( .ip1(n11855), .ip2(\cache_data_A[2][52] ), .op(n11621) );
  and2_1 U14551 ( .ip1(n12581), .ip2(\cache_data_A[7][52] ), .op(n11618) );
  nand2_1 U14552 ( .ip1(n11304), .ip2(\cache_data_A[5][52] ), .op(n11616) );
  nand2_1 U14553 ( .ip1(n12584), .ip2(\cache_data_A[4][52] ), .op(n11615) );
  nand2_1 U14554 ( .ip1(n11780), .ip2(\cache_data_A[6][52] ), .op(n11614) );
  nand2_1 U14555 ( .ip1(n12410), .ip2(\cache_data_A[3][52] ), .op(n11613) );
  nand4_1 U14556 ( .ip1(n11616), .ip2(n11615), .ip3(n11614), .ip4(n11613), 
        .op(n11617) );
  not_ab_or_c_or_d U14557 ( .ip1(\cache_data_A[0][52] ), .ip2(n12297), .ip3(
        n11618), .ip4(n11617), .op(n11620) );
  nand2_1 U14558 ( .ip1(n12242), .ip2(\cache_data_A[1][52] ), .op(n11619) );
  nand3_1 U14559 ( .ip1(n11621), .ip2(n11620), .ip3(n11619), .op(n12965) );
  nand2_1 U14560 ( .ip1(n12595), .ip2(n12965), .op(n11622) );
  nand4_1 U14561 ( .ip1(n11625), .ip2(n11624), .ip3(n11623), .ip4(n11622), 
        .op(n11626) );
  not_ab_or_c_or_d U14562 ( .ip1(n12563), .ip2(n12964), .ip3(n11627), .ip4(
        n11626), .op(n11638) );
  nand2_1 U14563 ( .ip1(\cache_data_B[2][20] ), .ip2(n12486), .op(n11636) );
  and2_1 U14564 ( .ip1(n12468), .ip2(\cache_data_B[7][20] ), .op(n11633) );
  nand2_1 U14565 ( .ip1(n12147), .ip2(\cache_data_B[1][20] ), .op(n11631) );
  nand2_1 U14566 ( .ip1(n12551), .ip2(\cache_data_B[6][20] ), .op(n11630) );
  nand2_1 U14567 ( .ip1(n12118), .ip2(\cache_data_B[5][20] ), .op(n11629) );
  nand2_1 U14568 ( .ip1(n12396), .ip2(\cache_data_B[4][20] ), .op(n11628) );
  nand4_1 U14569 ( .ip1(n11631), .ip2(n11630), .ip3(n11629), .ip4(n11628), 
        .op(n11632) );
  not_ab_or_c_or_d U14570 ( .ip1(\cache_data_B[0][20] ), .ip2(n12297), .ip3(
        n11633), .ip4(n11632), .op(n11635) );
  nand2_1 U14571 ( .ip1(n8060), .ip2(\cache_data_B[3][20] ), .op(n11634) );
  nand3_1 U14572 ( .ip1(n11636), .ip2(n11635), .ip3(n11634), .op(n12967) );
  nand2_1 U14573 ( .ip1(n12539), .ip2(n12967), .op(n11637) );
  nand3_1 U14574 ( .ip1(n11639), .ip2(n11638), .ip3(n11637), .op(n11640) );
  mux2_1 U14575 ( .ip1(N4144), .ip2(n11640), .s(n12599), .op(n5300) );
  nand2_1 U14576 ( .ip1(n12468), .ip2(\cache_data_A[7][53] ), .op(n11649) );
  and2_1 U14577 ( .ip1(n11156), .ip2(\cache_data_A[4][53] ), .op(n11646) );
  nand2_1 U14578 ( .ip1(n11780), .ip2(\cache_data_A[6][53] ), .op(n11644) );
  nand2_1 U14579 ( .ip1(n11855), .ip2(\cache_data_A[2][53] ), .op(n11643) );
  nand2_1 U14580 ( .ip1(n12147), .ip2(\cache_data_A[1][53] ), .op(n11642) );
  nand2_1 U14581 ( .ip1(n12591), .ip2(\cache_data_A[3][53] ), .op(n11641) );
  nand4_1 U14582 ( .ip1(n11644), .ip2(n11643), .ip3(n11642), .ip4(n11641), 
        .op(n11645) );
  not_ab_or_c_or_d U14583 ( .ip1(n12297), .ip2(\cache_data_A[0][53] ), .ip3(
        n11646), .ip4(n11645), .op(n11648) );
  nand2_1 U14584 ( .ip1(n12118), .ip2(\cache_data_A[5][53] ), .op(n11647) );
  nand3_1 U14585 ( .ip1(n11649), .ip2(n11648), .ip3(n11647), .op(n12992) );
  nand2_1 U14586 ( .ip1(n12595), .ip2(n12992), .op(n11722) );
  nand2_1 U14587 ( .ip1(n11911), .ip2(\cache_data_B[0][117] ), .op(n11658) );
  and2_1 U14588 ( .ip1(n12396), .ip2(\cache_data_B[4][117] ), .op(n11655) );
  nand2_1 U14589 ( .ip1(n12147), .ip2(\cache_data_B[1][117] ), .op(n11653) );
  nand2_1 U14590 ( .ip1(n11057), .ip2(\cache_data_B[7][117] ), .op(n11652) );
  nand2_1 U14591 ( .ip1(n11780), .ip2(\cache_data_B[6][117] ), .op(n11651) );
  nand2_1 U14592 ( .ip1(n12118), .ip2(\cache_data_B[5][117] ), .op(n11650) );
  nand4_1 U14593 ( .ip1(n11653), .ip2(n11652), .ip3(n11651), .ip4(n11650), 
        .op(n11654) );
  not_ab_or_c_or_d U14594 ( .ip1(n12546), .ip2(\cache_data_B[2][117] ), .ip3(
        n11655), .ip4(n11654), .op(n11657) );
  nand2_1 U14595 ( .ip1(n12321), .ip2(\cache_data_B[3][117] ), .op(n11656) );
  nand3_1 U14596 ( .ip1(n11658), .ip2(n11657), .ip3(n11656), .op(n12985) );
  nand2_1 U14597 ( .ip1(n12118), .ip2(\cache_data_A[5][85] ), .op(n11662) );
  nand2_1 U14598 ( .ip1(n12410), .ip2(\cache_data_A[3][85] ), .op(n11661) );
  nand2_1 U14599 ( .ip1(n12147), .ip2(\cache_data_A[1][85] ), .op(n11660) );
  nand2_1 U14600 ( .ip1(n12476), .ip2(\cache_data_A[4][85] ), .op(n11659) );
  nand4_1 U14601 ( .ip1(n11662), .ip2(n11661), .ip3(n11660), .ip4(n11659), 
        .op(n11668) );
  nand2_1 U14602 ( .ip1(n12581), .ip2(\cache_data_A[7][85] ), .op(n11666) );
  nand2_1 U14603 ( .ip1(n11780), .ip2(\cache_data_A[6][85] ), .op(n11665) );
  nand2_1 U14604 ( .ip1(n11855), .ip2(\cache_data_A[2][85] ), .op(n11664) );
  nand2_1 U14605 ( .ip1(n11911), .ip2(\cache_data_A[0][85] ), .op(n11663) );
  nand4_1 U14606 ( .ip1(n11666), .ip2(n11665), .ip3(n11664), .ip4(n11663), 
        .op(n11667) );
  nor2_1 U14607 ( .ip1(n11668), .ip2(n11667), .op(n12981) );
  nor2_1 U14608 ( .ip1(n12981), .ip2(n12529), .op(n11710) );
  nand2_1 U14609 ( .ip1(n11911), .ip2(\cache_data_B[0][21] ), .op(n11677) );
  and2_1 U14610 ( .ip1(n12256), .ip2(\cache_data_B[5][21] ), .op(n11674) );
  nand2_1 U14611 ( .ip1(n12054), .ip2(\cache_data_B[4][21] ), .op(n11672) );
  nand2_1 U14612 ( .ip1(n12321), .ip2(\cache_data_B[3][21] ), .op(n11671) );
  nand2_1 U14613 ( .ip1(n11855), .ip2(\cache_data_B[2][21] ), .op(n11670) );
  nand2_1 U14614 ( .ip1(n12429), .ip2(\cache_data_B[6][21] ), .op(n11669) );
  nand4_1 U14615 ( .ip1(n11672), .ip2(n11671), .ip3(n11670), .ip4(n11669), 
        .op(n11673) );
  not_ab_or_c_or_d U14616 ( .ip1(\cache_data_B[7][21] ), .ip2(n12278), .ip3(
        n11674), .ip4(n11673), .op(n11676) );
  nand2_1 U14617 ( .ip1(n12242), .ip2(\cache_data_B[1][21] ), .op(n11675) );
  nand3_1 U14618 ( .ip1(n11677), .ip2(n11676), .ip3(n11675), .op(n12980) );
  nand2_1 U14619 ( .ip1(n12539), .ip2(n12980), .op(n11708) );
  nand2_1 U14620 ( .ip1(n12147), .ip2(\cache_data_B[1][85] ), .op(n11686) );
  and2_1 U14621 ( .ip1(n12410), .ip2(\cache_data_B[3][85] ), .op(n11683) );
  nand2_1 U14622 ( .ip1(n11911), .ip2(\cache_data_B[0][85] ), .op(n11681) );
  nand2_1 U14623 ( .ip1(n10575), .ip2(\cache_data_B[7][85] ), .op(n11680) );
  nand2_1 U14624 ( .ip1(n11780), .ip2(\cache_data_B[6][85] ), .op(n11679) );
  nand2_1 U14625 ( .ip1(n11324), .ip2(\cache_data_B[4][85] ), .op(n11678) );
  nand4_1 U14626 ( .ip1(n11681), .ip2(n11680), .ip3(n11679), .ip4(n11678), 
        .op(n11682) );
  not_ab_or_c_or_d U14627 ( .ip1(\cache_data_B[2][85] ), .ip2(n12546), .ip3(
        n11683), .ip4(n11682), .op(n11685) );
  nand2_1 U14628 ( .ip1(n12256), .ip2(\cache_data_B[5][85] ), .op(n11684) );
  nand3_1 U14629 ( .ip1(n11686), .ip2(n11685), .ip3(n11684), .op(n12984) );
  nand2_1 U14630 ( .ip1(n12580), .ip2(n12984), .op(n11707) );
  nand2_1 U14631 ( .ip1(n11911), .ip2(\cache_data_A[0][21] ), .op(n11695) );
  and2_1 U14632 ( .ip1(n12256), .ip2(\cache_data_A[5][21] ), .op(n11692) );
  nand2_1 U14633 ( .ip1(n12321), .ip2(\cache_data_A[3][21] ), .op(n11690) );
  nand2_1 U14634 ( .ip1(n12371), .ip2(\cache_data_A[6][21] ), .op(n11689) );
  nand2_1 U14635 ( .ip1(n11855), .ip2(\cache_data_A[2][21] ), .op(n11688) );
  nand2_1 U14636 ( .ip1(n12476), .ip2(\cache_data_A[4][21] ), .op(n11687) );
  nand4_1 U14637 ( .ip1(n11690), .ip2(n11689), .ip3(n11688), .ip4(n11687), 
        .op(n11691) );
  not_ab_or_c_or_d U14638 ( .ip1(\cache_data_A[7][21] ), .ip2(n12278), .ip3(
        n11692), .ip4(n11691), .op(n11694) );
  nand2_1 U14639 ( .ip1(n12242), .ip2(\cache_data_A[1][21] ), .op(n11693) );
  nand3_1 U14640 ( .ip1(n11695), .ip2(n11694), .ip3(n11693), .op(n12982) );
  nand2_1 U14641 ( .ip1(n12550), .ip2(n12982), .op(n11706) );
  nand2_1 U14642 ( .ip1(n12581), .ip2(\cache_data_A[7][117] ), .op(n11704) );
  and2_1 U14643 ( .ip1(n11946), .ip2(\cache_data_A[1][117] ), .op(n11701) );
  nand2_1 U14644 ( .ip1(n12118), .ip2(\cache_data_A[5][117] ), .op(n11699) );
  nand2_1 U14645 ( .ip1(n11855), .ip2(\cache_data_A[2][117] ), .op(n11698) );
  nand2_1 U14646 ( .ip1(n12194), .ip2(\cache_data_A[4][117] ), .op(n11697) );
  nand2_1 U14647 ( .ip1(n11911), .ip2(\cache_data_A[0][117] ), .op(n11696) );
  nand4_1 U14648 ( .ip1(n11699), .ip2(n11698), .ip3(n11697), .ip4(n11696), 
        .op(n11700) );
  not_ab_or_c_or_d U14649 ( .ip1(\cache_data_A[6][117] ), .ip2(n12337), .ip3(
        n11701), .ip4(n11700), .op(n11703) );
  nand2_1 U14650 ( .ip1(n12321), .ip2(\cache_data_A[3][117] ), .op(n11702) );
  nand3_1 U14651 ( .ip1(n11704), .ip2(n11703), .ip3(n11702), .op(n12983) );
  nand2_1 U14652 ( .ip1(n12509), .ip2(n12983), .op(n11705) );
  nand4_1 U14653 ( .ip1(n11708), .ip2(n11707), .ip3(n11706), .ip4(n11705), 
        .op(n11709) );
  not_ab_or_c_or_d U14654 ( .ip1(n12573), .ip2(n12985), .ip3(n11710), .ip4(
        n11709), .op(n11721) );
  nand2_1 U14655 ( .ip1(n12429), .ip2(\cache_data_B[6][53] ), .op(n11719) );
  and2_1 U14656 ( .ip1(n12486), .ip2(\cache_data_B[2][53] ), .op(n11716) );
  nand2_1 U14657 ( .ip1(n11280), .ip2(\cache_data_B[5][53] ), .op(n11714) );
  nand2_1 U14658 ( .ip1(n8060), .ip2(\cache_data_B[3][53] ), .op(n11713) );
  nand2_1 U14659 ( .ip1(n12581), .ip2(\cache_data_B[7][53] ), .op(n11712) );
  nand2_1 U14660 ( .ip1(n12147), .ip2(\cache_data_B[1][53] ), .op(n11711) );
  nand4_1 U14661 ( .ip1(n11714), .ip2(n11713), .ip3(n11712), .ip4(n11711), 
        .op(n11715) );
  not_ab_or_c_or_d U14662 ( .ip1(\cache_data_B[0][53] ), .ip2(n12297), .ip3(
        n11716), .ip4(n11715), .op(n11718) );
  nand2_1 U14663 ( .ip1(n12194), .ip2(\cache_data_B[4][53] ), .op(n11717) );
  nand3_1 U14664 ( .ip1(n11719), .ip2(n11718), .ip3(n11717), .op(n12993) );
  nand2_1 U14665 ( .ip1(n12563), .ip2(n12993), .op(n11720) );
  nand3_1 U14666 ( .ip1(n11722), .ip2(n11721), .ip3(n11720), .op(n11723) );
  mux2_1 U14667 ( .ip1(N4141), .ip2(n11723), .s(n12599), .op(n5299) );
  nand2_1 U14668 ( .ip1(n11780), .ip2(\cache_data_A[6][118] ), .op(n11733) );
  and2_1 U14669 ( .ip1(n12468), .ip2(\cache_data_A[7][118] ), .op(n11730) );
  nand2_1 U14670 ( .ip1(n11855), .ip2(\cache_data_A[2][118] ), .op(n11728) );
  nand2_1 U14671 ( .ip1(n11724), .ip2(\cache_data_A[1][118] ), .op(n11727) );
  nand2_1 U14672 ( .ip1(n11304), .ip2(\cache_data_A[5][118] ), .op(n11726) );
  nand2_1 U14673 ( .ip1(n12396), .ip2(\cache_data_A[4][118] ), .op(n11725) );
  nand4_1 U14674 ( .ip1(n11728), .ip2(n11727), .ip3(n11726), .ip4(n11725), 
        .op(n11729) );
  not_ab_or_c_or_d U14675 ( .ip1(\cache_data_A[0][118] ), .ip2(n12297), .ip3(
        n11730), .ip4(n11729), .op(n11732) );
  nand2_1 U14676 ( .ip1(n12321), .ip2(\cache_data_A[3][118] ), .op(n11731) );
  nand3_1 U14677 ( .ip1(n11733), .ip2(n11732), .ip3(n11731), .op(n13000) );
  nand2_1 U14678 ( .ip1(n12509), .ip2(n13000), .op(n11807) );
  nand2_1 U14679 ( .ip1(n12429), .ip2(\cache_data_A[6][22] ), .op(n11742) );
  and2_1 U14680 ( .ip1(n12410), .ip2(\cache_data_A[3][22] ), .op(n11739) );
  nand2_1 U14681 ( .ip1(n11855), .ip2(\cache_data_A[2][22] ), .op(n11737) );
  nand2_1 U14682 ( .ip1(n11156), .ip2(\cache_data_A[4][22] ), .op(n11736) );
  nand2_1 U14683 ( .ip1(n11911), .ip2(\cache_data_A[0][22] ), .op(n11735) );
  nand2_1 U14684 ( .ip1(n12256), .ip2(\cache_data_A[5][22] ), .op(n11734) );
  nand4_1 U14685 ( .ip1(n11737), .ip2(n11736), .ip3(n11735), .ip4(n11734), 
        .op(n11738) );
  not_ab_or_c_or_d U14686 ( .ip1(\cache_data_A[7][22] ), .ip2(n11057), .ip3(
        n11739), .ip4(n11738), .op(n11741) );
  nand2_1 U14687 ( .ip1(n12242), .ip2(\cache_data_A[1][22] ), .op(n11740) );
  nand3_1 U14688 ( .ip1(n11742), .ip2(n11741), .ip3(n11740), .op(n13001) );
  nand2_1 U14689 ( .ip1(n12118), .ip2(\cache_data_A[5][86] ), .op(n11746) );
  nand2_1 U14690 ( .ip1(n11911), .ip2(\cache_data_A[0][86] ), .op(n11745) );
  nand2_1 U14691 ( .ip1(n12429), .ip2(\cache_data_A[6][86] ), .op(n11744) );
  nand2_1 U14692 ( .ip1(n12194), .ip2(\cache_data_A[4][86] ), .op(n11743) );
  nand4_1 U14693 ( .ip1(n11746), .ip2(n11745), .ip3(n11744), .ip4(n11743), 
        .op(n11752) );
  nand2_1 U14694 ( .ip1(n12147), .ip2(\cache_data_A[1][86] ), .op(n11750) );
  nand2_1 U14695 ( .ip1(n12581), .ip2(\cache_data_A[7][86] ), .op(n11749) );
  nand2_1 U14696 ( .ip1(n11855), .ip2(\cache_data_A[2][86] ), .op(n11748) );
  nand2_1 U14697 ( .ip1(n8060), .ip2(\cache_data_A[3][86] ), .op(n11747) );
  nand4_1 U14698 ( .ip1(n11750), .ip2(n11749), .ip3(n11748), .ip4(n11747), 
        .op(n11751) );
  nor2_1 U14699 ( .ip1(n11752), .ip2(n11751), .op(n12999) );
  nor2_1 U14700 ( .ip1(n12999), .ip2(n12529), .op(n11795) );
  nand2_1 U14701 ( .ip1(n12321), .ip2(\cache_data_B[3][118] ), .op(n11761) );
  and2_1 U14702 ( .ip1(n10686), .ip2(\cache_data_B[1][118] ), .op(n11758) );
  nand2_1 U14703 ( .ip1(n12194), .ip2(\cache_data_B[4][118] ), .op(n11756) );
  nand2_1 U14704 ( .ip1(n11911), .ip2(\cache_data_B[0][118] ), .op(n11755) );
  nand2_1 U14705 ( .ip1(n10575), .ip2(\cache_data_B[7][118] ), .op(n11754) );
  nand2_1 U14706 ( .ip1(n12371), .ip2(\cache_data_B[6][118] ), .op(n11753) );
  nand4_1 U14707 ( .ip1(n11756), .ip2(n11755), .ip3(n11754), .ip4(n11753), 
        .op(n11757) );
  not_ab_or_c_or_d U14708 ( .ip1(n12475), .ip2(\cache_data_B[2][118] ), .ip3(
        n11758), .ip4(n11757), .op(n11760) );
  nand2_1 U14709 ( .ip1(n12118), .ip2(\cache_data_B[5][118] ), .op(n11759) );
  nand3_1 U14710 ( .ip1(n11761), .ip2(n11760), .ip3(n11759), .op(n13002) );
  nand2_1 U14711 ( .ip1(n12573), .ip2(n13002), .op(n11793) );
  nand2_1 U14712 ( .ip1(n11855), .ip2(\cache_data_B[2][22] ), .op(n11770) );
  and2_1 U14713 ( .ip1(n12582), .ip2(\cache_data_B[5][22] ), .op(n11767) );
  nand2_1 U14714 ( .ip1(n12410), .ip2(\cache_data_B[3][22] ), .op(n11765) );
  nand2_1 U14715 ( .ip1(n11911), .ip2(\cache_data_B[0][22] ), .op(n11764) );
  nand2_1 U14716 ( .ip1(n10702), .ip2(\cache_data_B[7][22] ), .op(n11763) );
  nand2_1 U14717 ( .ip1(n12147), .ip2(\cache_data_B[1][22] ), .op(n11762) );
  nand4_1 U14718 ( .ip1(n11765), .ip2(n11764), .ip3(n11763), .ip4(n11762), 
        .op(n11766) );
  not_ab_or_c_or_d U14719 ( .ip1(\cache_data_B[6][22] ), .ip2(n12320), .ip3(
        n11767), .ip4(n11766), .op(n11769) );
  nand2_1 U14720 ( .ip1(n12476), .ip2(\cache_data_B[4][22] ), .op(n11768) );
  nand3_1 U14721 ( .ip1(n11770), .ip2(n11769), .ip3(n11768), .op(n13003) );
  nand2_1 U14722 ( .ip1(n12539), .ip2(n13003), .op(n11792) );
  nand2_1 U14723 ( .ip1(n12321), .ip2(\cache_data_B[3][86] ), .op(n11779) );
  and2_1 U14724 ( .ip1(n12147), .ip2(\cache_data_B[1][86] ), .op(n11776) );
  nand2_1 U14725 ( .ip1(n12582), .ip2(\cache_data_B[5][86] ), .op(n11774) );
  nand2_1 U14726 ( .ip1(n11911), .ip2(\cache_data_B[0][86] ), .op(n11773) );
  nand2_1 U14727 ( .ip1(n10575), .ip2(\cache_data_B[7][86] ), .op(n11772) );
  nand2_1 U14728 ( .ip1(n11855), .ip2(\cache_data_B[2][86] ), .op(n11771) );
  nand4_1 U14729 ( .ip1(n11774), .ip2(n11773), .ip3(n11772), .ip4(n11771), 
        .op(n11775) );
  not_ab_or_c_or_d U14730 ( .ip1(\cache_data_B[6][86] ), .ip2(n12337), .ip3(
        n11776), .ip4(n11775), .op(n11778) );
  nand2_1 U14731 ( .ip1(n12194), .ip2(\cache_data_B[4][86] ), .op(n11777) );
  nand3_1 U14732 ( .ip1(n11779), .ip2(n11778), .ip3(n11777), .op(n12998) );
  nand2_1 U14733 ( .ip1(n12580), .ip2(n12998), .op(n11791) );
  nand2_1 U14734 ( .ip1(n11855), .ip2(\cache_data_B[2][54] ), .op(n11789) );
  and2_1 U14735 ( .ip1(n11280), .ip2(\cache_data_B[5][54] ), .op(n11786) );
  nand2_1 U14736 ( .ip1(n11911), .ip2(\cache_data_B[0][54] ), .op(n11784) );
  nand2_1 U14737 ( .ip1(n11780), .ip2(\cache_data_B[6][54] ), .op(n11783) );
  nand2_1 U14738 ( .ip1(n11324), .ip2(\cache_data_B[4][54] ), .op(n11782) );
  nand2_1 U14739 ( .ip1(n10575), .ip2(\cache_data_B[7][54] ), .op(n11781) );
  nand4_1 U14740 ( .ip1(n11784), .ip2(n11783), .ip3(n11782), .ip4(n11781), 
        .op(n11785) );
  not_ab_or_c_or_d U14741 ( .ip1(n12096), .ip2(\cache_data_B[3][54] ), .ip3(
        n11786), .ip4(n11785), .op(n11788) );
  nand2_1 U14742 ( .ip1(n12242), .ip2(\cache_data_B[1][54] ), .op(n11787) );
  nand3_1 U14743 ( .ip1(n11789), .ip2(n11788), .ip3(n11787), .op(n13010) );
  nand2_1 U14744 ( .ip1(n12563), .ip2(n13010), .op(n11790) );
  nand4_1 U14745 ( .ip1(n11793), .ip2(n11792), .ip3(n11791), .ip4(n11790), 
        .op(n11794) );
  not_ab_or_c_or_d U14746 ( .ip1(n12550), .ip2(n13001), .ip3(n11795), .ip4(
        n11794), .op(n11806) );
  nand2_1 U14747 ( .ip1(n12429), .ip2(\cache_data_A[6][54] ), .op(n11804) );
  and2_1 U14748 ( .ip1(n12321), .ip2(\cache_data_A[3][54] ), .op(n11801) );
  nand2_1 U14749 ( .ip1(n12581), .ip2(\cache_data_A[7][54] ), .op(n11799) );
  nand2_1 U14750 ( .ip1(n11855), .ip2(\cache_data_A[2][54] ), .op(n11798) );
  nand2_1 U14751 ( .ip1(n11296), .ip2(\cache_data_A[5][54] ), .op(n11797) );
  nand2_1 U14752 ( .ip1(n12242), .ip2(\cache_data_A[1][54] ), .op(n11796) );
  nand4_1 U14753 ( .ip1(n11799), .ip2(n11798), .ip3(n11797), .ip4(n11796), 
        .op(n11800) );
  not_ab_or_c_or_d U14754 ( .ip1(\cache_data_A[0][54] ), .ip2(n8452), .ip3(
        n11801), .ip4(n11800), .op(n11803) );
  nand2_1 U14755 ( .ip1(n12476), .ip2(\cache_data_A[4][54] ), .op(n11802) );
  nand3_1 U14756 ( .ip1(n11804), .ip2(n11803), .ip3(n11802), .op(n13011) );
  nand2_1 U14757 ( .ip1(n12595), .ip2(n13011), .op(n11805) );
  nand3_1 U14758 ( .ip1(n11807), .ip2(n11806), .ip3(n11805), .op(n11808) );
  mux2_1 U14759 ( .ip1(N4138), .ip2(n11808), .s(n12599), .op(n5298) );
  nand2_1 U14760 ( .ip1(n11911), .ip2(\cache_data_A[0][119] ), .op(n11817) );
  and2_1 U14761 ( .ip1(n11296), .ip2(\cache_data_A[5][119] ), .op(n11814) );
  nand2_1 U14762 ( .ip1(n12321), .ip2(\cache_data_A[3][119] ), .op(n11812) );
  nand2_1 U14763 ( .ip1(n12429), .ip2(\cache_data_A[6][119] ), .op(n11811) );
  nand2_1 U14764 ( .ip1(n11855), .ip2(\cache_data_A[2][119] ), .op(n11810) );
  nand2_1 U14765 ( .ip1(n12476), .ip2(\cache_data_A[4][119] ), .op(n11809) );
  nand4_1 U14766 ( .ip1(n11812), .ip2(n11811), .ip3(n11810), .ip4(n11809), 
        .op(n11813) );
  not_ab_or_c_or_d U14767 ( .ip1(\cache_data_A[1][119] ), .ip2(n11946), .ip3(
        n11814), .ip4(n11813), .op(n11816) );
  nand2_1 U14768 ( .ip1(n12468), .ip2(\cache_data_A[7][119] ), .op(n11815) );
  nand3_1 U14769 ( .ip1(n11817), .ip2(n11816), .ip3(n11815), .op(n13016) );
  nand2_1 U14770 ( .ip1(n12509), .ip2(n13016), .op(n11891) );
  nand2_1 U14771 ( .ip1(n11911), .ip2(\cache_data_B[0][87] ), .op(n11826) );
  and2_1 U14772 ( .ip1(n12194), .ip2(\cache_data_B[4][87] ), .op(n11823) );
  nand2_1 U14773 ( .ip1(n10702), .ip2(\cache_data_B[7][87] ), .op(n11821) );
  nand2_1 U14774 ( .ip1(n12321), .ip2(\cache_data_B[3][87] ), .op(n11820) );
  nand2_1 U14775 ( .ip1(n12242), .ip2(\cache_data_B[1][87] ), .op(n11819) );
  nand2_1 U14776 ( .ip1(n11280), .ip2(\cache_data_B[5][87] ), .op(n11818) );
  nand4_1 U14777 ( .ip1(n11821), .ip2(n11820), .ip3(n11819), .ip4(n11818), 
        .op(n11822) );
  not_ab_or_c_or_d U14778 ( .ip1(\cache_data_B[2][87] ), .ip2(n12546), .ip3(
        n11823), .ip4(n11822), .op(n11825) );
  nand2_1 U14779 ( .ip1(n12429), .ip2(\cache_data_B[6][87] ), .op(n11824) );
  nand3_1 U14780 ( .ip1(n11826), .ip2(n11825), .ip3(n11824), .op(n13029) );
  nand2_1 U14781 ( .ip1(n12429), .ip2(\cache_data_A[6][87] ), .op(n11830) );
  nand2_1 U14782 ( .ip1(n11855), .ip2(\cache_data_A[2][87] ), .op(n11829) );
  nand2_1 U14783 ( .ip1(n12410), .ip2(\cache_data_A[3][87] ), .op(n11828) );
  nand2_1 U14784 ( .ip1(n12476), .ip2(\cache_data_A[4][87] ), .op(n11827) );
  nand4_1 U14785 ( .ip1(n11830), .ip2(n11829), .ip3(n11828), .ip4(n11827), 
        .op(n11836) );
  nand2_1 U14786 ( .ip1(n12242), .ip2(\cache_data_A[1][87] ), .op(n11834) );
  nand2_1 U14787 ( .ip1(n11911), .ip2(\cache_data_A[0][87] ), .op(n11833) );
  nand2_1 U14788 ( .ip1(n10702), .ip2(\cache_data_A[7][87] ), .op(n11832) );
  nand2_1 U14789 ( .ip1(n12256), .ip2(\cache_data_A[5][87] ), .op(n11831) );
  nand4_1 U14790 ( .ip1(n11834), .ip2(n11833), .ip3(n11832), .ip4(n11831), 
        .op(n11835) );
  nor2_1 U14791 ( .ip1(n11836), .ip2(n11835), .op(n13017) );
  nor2_1 U14792 ( .ip1(n13017), .ip2(n12529), .op(n11879) );
  nand2_1 U14793 ( .ip1(n12429), .ip2(\cache_data_A[6][23] ), .op(n11845) );
  and2_1 U14794 ( .ip1(n11946), .ip2(\cache_data_A[1][23] ), .op(n11842) );
  nand2_1 U14795 ( .ip1(n11911), .ip2(\cache_data_A[0][23] ), .op(n11840) );
  nand2_1 U14796 ( .ip1(n10575), .ip2(\cache_data_A[7][23] ), .op(n11839) );
  nand2_1 U14797 ( .ip1(n11855), .ip2(\cache_data_A[2][23] ), .op(n11838) );
  nand2_1 U14798 ( .ip1(n8060), .ip2(\cache_data_A[3][23] ), .op(n11837) );
  nand4_1 U14799 ( .ip1(n11840), .ip2(n11839), .ip3(n11838), .ip4(n11837), 
        .op(n11841) );
  not_ab_or_c_or_d U14800 ( .ip1(n12396), .ip2(\cache_data_A[4][23] ), .ip3(
        n11842), .ip4(n11841), .op(n11844) );
  nand2_1 U14801 ( .ip1(n11296), .ip2(\cache_data_A[5][23] ), .op(n11843) );
  nand3_1 U14802 ( .ip1(n11845), .ip2(n11844), .ip3(n11843), .op(n13019) );
  nand2_1 U14803 ( .ip1(n12550), .ip2(n13019), .op(n11877) );
  nand2_1 U14804 ( .ip1(n10702), .ip2(\cache_data_B[7][23] ), .op(n11854) );
  and2_1 U14805 ( .ip1(n12591), .ip2(\cache_data_B[3][23] ), .op(n11851) );
  nand2_1 U14806 ( .ip1(n11296), .ip2(\cache_data_B[5][23] ), .op(n11849) );
  nand2_1 U14807 ( .ip1(n12429), .ip2(\cache_data_B[6][23] ), .op(n11848) );
  nand2_1 U14808 ( .ip1(n11855), .ip2(\cache_data_B[2][23] ), .op(n11847) );
  nand2_1 U14809 ( .ip1(n12396), .ip2(\cache_data_B[4][23] ), .op(n11846) );
  nand4_1 U14810 ( .ip1(n11849), .ip2(n11848), .ip3(n11847), .ip4(n11846), 
        .op(n11850) );
  not_ab_or_c_or_d U14811 ( .ip1(\cache_data_B[0][23] ), .ip2(n8452), .ip3(
        n11851), .ip4(n11850), .op(n11853) );
  nand2_1 U14812 ( .ip1(n12242), .ip2(\cache_data_B[1][23] ), .op(n11852) );
  nand3_1 U14813 ( .ip1(n11854), .ip2(n11853), .ip3(n11852), .op(n13028) );
  nand2_1 U14814 ( .ip1(n12539), .ip2(n13028), .op(n11876) );
  nand2_1 U14815 ( .ip1(n11057), .ip2(\cache_data_B[7][55] ), .op(n11864) );
  and2_1 U14816 ( .ip1(n12194), .ip2(\cache_data_B[4][55] ), .op(n11861) );
  nand2_1 U14817 ( .ip1(n11304), .ip2(\cache_data_B[5][55] ), .op(n11859) );
  nand2_1 U14818 ( .ip1(n12242), .ip2(\cache_data_B[1][55] ), .op(n11858) );
  nand2_1 U14819 ( .ip1(n11911), .ip2(\cache_data_B[0][55] ), .op(n11857) );
  nand2_1 U14820 ( .ip1(n11855), .ip2(\cache_data_B[2][55] ), .op(n11856) );
  nand4_1 U14821 ( .ip1(n11859), .ip2(n11858), .ip3(n11857), .ip4(n11856), 
        .op(n11860) );
  not_ab_or_c_or_d U14822 ( .ip1(n12096), .ip2(\cache_data_B[3][55] ), .ip3(
        n11861), .ip4(n11860), .op(n11863) );
  nand2_1 U14823 ( .ip1(n12429), .ip2(\cache_data_B[6][55] ), .op(n11862) );
  nand3_1 U14824 ( .ip1(n11864), .ip2(n11863), .ip3(n11862), .op(n13020) );
  nand2_1 U14825 ( .ip1(n12563), .ip2(n13020), .op(n11875) );
  nand2_1 U14826 ( .ip1(\cache_data_A[2][55] ), .ip2(n12486), .op(n11873) );
  and2_1 U14827 ( .ip1(n11296), .ip2(\cache_data_A[5][55] ), .op(n11870) );
  nand2_1 U14828 ( .ip1(n12242), .ip2(\cache_data_A[1][55] ), .op(n11868) );
  nand2_1 U14829 ( .ip1(n11057), .ip2(\cache_data_A[7][55] ), .op(n11867) );
  nand2_1 U14830 ( .ip1(n11911), .ip2(\cache_data_A[0][55] ), .op(n11866) );
  nand2_1 U14831 ( .ip1(n8060), .ip2(\cache_data_A[3][55] ), .op(n11865) );
  nand4_1 U14832 ( .ip1(n11868), .ip2(n11867), .ip3(n11866), .ip4(n11865), 
        .op(n11869) );
  not_ab_or_c_or_d U14833 ( .ip1(n12551), .ip2(\cache_data_A[6][55] ), .ip3(
        n11870), .ip4(n11869), .op(n11872) );
  nand2_1 U14834 ( .ip1(n12476), .ip2(\cache_data_A[4][55] ), .op(n11871) );
  nand3_1 U14835 ( .ip1(n11873), .ip2(n11872), .ip3(n11871), .op(n13018) );
  nand2_1 U14836 ( .ip1(n12595), .ip2(n13018), .op(n11874) );
  nand4_1 U14837 ( .ip1(n11877), .ip2(n11876), .ip3(n11875), .ip4(n11874), 
        .op(n11878) );
  not_ab_or_c_or_d U14838 ( .ip1(n12580), .ip2(n13029), .ip3(n11879), .ip4(
        n11878), .op(n11890) );
  nand2_1 U14839 ( .ip1(\cache_data_B[4][119] ), .ip2(n12584), .op(n11888) );
  and2_1 U14840 ( .ip1(n12429), .ip2(\cache_data_B[6][119] ), .op(n11885) );
  nand2_1 U14841 ( .ip1(n12559), .ip2(\cache_data_B[3][119] ), .op(n11883) );
  nand2_1 U14842 ( .ip1(n10575), .ip2(\cache_data_B[7][119] ), .op(n11882) );
  nand2_1 U14843 ( .ip1(n12475), .ip2(\cache_data_B[2][119] ), .op(n11881) );
  nand2_1 U14844 ( .ip1(n12242), .ip2(\cache_data_B[1][119] ), .op(n11880) );
  nand4_1 U14845 ( .ip1(n11883), .ip2(n11882), .ip3(n11881), .ip4(n11880), 
        .op(n11884) );
  not_ab_or_c_or_d U14846 ( .ip1(n12297), .ip2(\cache_data_B[0][119] ), .ip3(
        n11885), .ip4(n11884), .op(n11887) );
  nand2_1 U14847 ( .ip1(n11296), .ip2(\cache_data_B[5][119] ), .op(n11886) );
  nand3_1 U14848 ( .ip1(n11888), .ip2(n11887), .ip3(n11886), .op(n13021) );
  nand2_1 U14849 ( .ip1(n12573), .ip2(n13021), .op(n11889) );
  nand3_1 U14850 ( .ip1(n11891), .ip2(n11890), .ip3(n11889), .op(n11892) );
  mux2_1 U14851 ( .ip1(N4135), .ip2(n11892), .s(n12599), .op(n5297) );
  nand2_1 U14852 ( .ip1(n12429), .ip2(\cache_data_B[6][88] ), .op(n11901) );
  and2_1 U14853 ( .ip1(n12118), .ip2(\cache_data_B[5][88] ), .op(n11898) );
  nand2_1 U14854 ( .ip1(n12242), .ip2(\cache_data_B[1][88] ), .op(n11896) );
  nand2_1 U14855 ( .ip1(n10575), .ip2(\cache_data_B[7][88] ), .op(n11895) );
  nand2_1 U14856 ( .ip1(n11855), .ip2(\cache_data_B[2][88] ), .op(n11894) );
  nand2_1 U14857 ( .ip1(n11911), .ip2(\cache_data_B[0][88] ), .op(n11893) );
  nand4_1 U14858 ( .ip1(n11896), .ip2(n11895), .ip3(n11894), .ip4(n11893), 
        .op(n11897) );
  not_ab_or_c_or_d U14859 ( .ip1(\cache_data_B[4][88] ), .ip2(n11156), .ip3(
        n11898), .ip4(n11897), .op(n11900) );
  nand2_1 U14860 ( .ip1(n12410), .ip2(\cache_data_B[3][88] ), .op(n11899) );
  nand3_1 U14861 ( .ip1(n11901), .ip2(n11900), .ip3(n11899), .op(n13048) );
  nand2_1 U14862 ( .ip1(n12580), .ip2(n13048), .op(n11976) );
  nand2_1 U14863 ( .ip1(n11057), .ip2(\cache_data_B[7][24] ), .op(n11910) );
  and2_1 U14864 ( .ip1(n12321), .ip2(\cache_data_B[3][24] ), .op(n11907) );
  nand2_1 U14865 ( .ip1(n11156), .ip2(\cache_data_B[4][24] ), .op(n11905) );
  nand2_1 U14866 ( .ip1(n12118), .ip2(\cache_data_B[5][24] ), .op(n11904) );
  nand2_1 U14867 ( .ip1(n12475), .ip2(\cache_data_B[2][24] ), .op(n11903) );
  nand2_1 U14868 ( .ip1(n12242), .ip2(\cache_data_B[1][24] ), .op(n11902) );
  nand4_1 U14869 ( .ip1(n11905), .ip2(n11904), .ip3(n11903), .ip4(n11902), 
        .op(n11906) );
  not_ab_or_c_or_d U14870 ( .ip1(\cache_data_B[0][24] ), .ip2(n12204), .ip3(
        n11907), .ip4(n11906), .op(n11909) );
  nand2_1 U14871 ( .ip1(n12429), .ip2(\cache_data_B[6][24] ), .op(n11908) );
  nand3_1 U14872 ( .ip1(n11910), .ip2(n11909), .ip3(n11908), .op(n13038) );
  nand2_1 U14873 ( .ip1(n12429), .ip2(\cache_data_A[6][88] ), .op(n11915) );
  nand2_1 U14874 ( .ip1(n12486), .ip2(\cache_data_A[2][88] ), .op(n11914) );
  nand2_1 U14875 ( .ip1(n12476), .ip2(\cache_data_A[4][88] ), .op(n11913) );
  nand2_1 U14876 ( .ip1(n11911), .ip2(\cache_data_A[0][88] ), .op(n11912) );
  nand4_1 U14877 ( .ip1(n11915), .ip2(n11914), .ip3(n11913), .ip4(n11912), 
        .op(n11921) );
  nand2_1 U14878 ( .ip1(n12410), .ip2(\cache_data_A[3][88] ), .op(n11919) );
  nand2_1 U14879 ( .ip1(n12468), .ip2(\cache_data_A[7][88] ), .op(n11918) );
  nand2_1 U14880 ( .ip1(n12242), .ip2(\cache_data_A[1][88] ), .op(n11917) );
  nand2_1 U14881 ( .ip1(n12582), .ip2(\cache_data_A[5][88] ), .op(n11916) );
  nand4_1 U14882 ( .ip1(n11919), .ip2(n11918), .ip3(n11917), .ip4(n11916), 
        .op(n11920) );
  nor2_1 U14883 ( .ip1(n11921), .ip2(n11920), .op(n13036) );
  nor2_1 U14884 ( .ip1(n13036), .ip2(n12529), .op(n11964) );
  nand2_1 U14885 ( .ip1(\cache_data_B[0][56] ), .ip2(n12204), .op(n11930) );
  and2_1 U14886 ( .ip1(n12147), .ip2(\cache_data_B[1][56] ), .op(n11927) );
  nand2_1 U14887 ( .ip1(n8060), .ip2(\cache_data_B[3][56] ), .op(n11925) );
  nand2_1 U14888 ( .ip1(n12582), .ip2(\cache_data_B[5][56] ), .op(n11924) );
  nand2_1 U14889 ( .ip1(n10702), .ip2(\cache_data_B[7][56] ), .op(n11923) );
  nand2_1 U14890 ( .ip1(n12396), .ip2(\cache_data_B[4][56] ), .op(n11922) );
  nand4_1 U14891 ( .ip1(n11925), .ip2(n11924), .ip3(n11923), .ip4(n11922), 
        .op(n11926) );
  not_ab_or_c_or_d U14892 ( .ip1(n12551), .ip2(\cache_data_B[6][56] ), .ip3(
        n11927), .ip4(n11926), .op(n11929) );
  nand2_1 U14893 ( .ip1(n11142), .ip2(\cache_data_B[2][56] ), .op(n11928) );
  nand3_1 U14894 ( .ip1(n11930), .ip2(n11929), .ip3(n11928), .op(n13039) );
  nand2_1 U14895 ( .ip1(n12563), .ip2(n13039), .op(n11962) );
  nand2_1 U14896 ( .ip1(\cache_data_B[6][120] ), .ip2(n12371), .op(n11939) );
  and2_1 U14897 ( .ip1(n12591), .ip2(\cache_data_B[3][120] ), .op(n11936) );
  nand2_1 U14898 ( .ip1(n12242), .ip2(\cache_data_B[1][120] ), .op(n11934) );
  nand2_1 U14899 ( .ip1(n12204), .ip2(\cache_data_B[0][120] ), .op(n11933) );
  nand2_1 U14900 ( .ip1(n11156), .ip2(\cache_data_B[4][120] ), .op(n11932) );
  nand2_1 U14901 ( .ip1(n12475), .ip2(\cache_data_B[2][120] ), .op(n11931) );
  nand4_1 U14902 ( .ip1(n11934), .ip2(n11933), .ip3(n11932), .ip4(n11931), 
        .op(n11935) );
  not_ab_or_c_or_d U14903 ( .ip1(\cache_data_B[7][120] ), .ip2(n10575), .ip3(
        n11936), .ip4(n11935), .op(n11938) );
  nand2_1 U14904 ( .ip1(n12582), .ip2(\cache_data_B[5][120] ), .op(n11937) );
  nand3_1 U14905 ( .ip1(n11939), .ip2(n11938), .ip3(n11937), .op(n13037) );
  nand2_1 U14906 ( .ip1(n12573), .ip2(n13037), .op(n11961) );
  nand2_1 U14907 ( .ip1(\cache_data_A[0][120] ), .ip2(n12204), .op(n11949) );
  and2_1 U14908 ( .ip1(n11296), .ip2(\cache_data_A[5][120] ), .op(n11945) );
  nand2_1 U14909 ( .ip1(n12429), .ip2(\cache_data_A[6][120] ), .op(n11943) );
  nand2_1 U14910 ( .ip1(n10575), .ip2(\cache_data_A[7][120] ), .op(n11942) );
  nand2_1 U14911 ( .ip1(n8060), .ip2(\cache_data_A[3][120] ), .op(n11941) );
  nand2_1 U14912 ( .ip1(n11324), .ip2(\cache_data_A[4][120] ), .op(n11940) );
  nand4_1 U14913 ( .ip1(n11943), .ip2(n11942), .ip3(n11941), .ip4(n11940), 
        .op(n11944) );
  not_ab_or_c_or_d U14914 ( .ip1(\cache_data_A[1][120] ), .ip2(n11946), .ip3(
        n11945), .ip4(n11944), .op(n11948) );
  nand2_1 U14915 ( .ip1(n11142), .ip2(\cache_data_A[2][120] ), .op(n11947) );
  nand3_1 U14916 ( .ip1(n11949), .ip2(n11948), .ip3(n11947), .op(n13040) );
  nand2_1 U14917 ( .ip1(n12509), .ip2(n13040), .op(n11960) );
  nand2_1 U14918 ( .ip1(n12242), .ip2(\cache_data_A[1][24] ), .op(n11958) );
  and2_1 U14919 ( .ip1(n12458), .ip2(\cache_data_A[6][24] ), .op(n11955) );
  nand2_1 U14920 ( .ip1(n11156), .ip2(\cache_data_A[4][24] ), .op(n11953) );
  nand2_1 U14921 ( .ip1(n12591), .ip2(\cache_data_A[3][24] ), .op(n11952) );
  nand2_1 U14922 ( .ip1(n12475), .ip2(\cache_data_A[2][24] ), .op(n11951) );
  nand2_1 U14923 ( .ip1(n12552), .ip2(\cache_data_A[7][24] ), .op(n11950) );
  nand4_1 U14924 ( .ip1(n11953), .ip2(n11952), .ip3(n11951), .ip4(n11950), 
        .op(n11954) );
  not_ab_or_c_or_d U14925 ( .ip1(n12297), .ip2(\cache_data_A[0][24] ), .ip3(
        n11955), .ip4(n11954), .op(n11957) );
  nand2_1 U14926 ( .ip1(n12582), .ip2(\cache_data_A[5][24] ), .op(n11956) );
  nand3_1 U14927 ( .ip1(n11958), .ip2(n11957), .ip3(n11956), .op(n13035) );
  nand2_1 U14928 ( .ip1(n12550), .ip2(n13035), .op(n11959) );
  nand4_1 U14929 ( .ip1(n11962), .ip2(n11961), .ip3(n11960), .ip4(n11959), 
        .op(n11963) );
  not_ab_or_c_or_d U14930 ( .ip1(n12539), .ip2(n13038), .ip3(n11964), .ip4(
        n11963), .op(n11975) );
  nand2_1 U14931 ( .ip1(\cache_data_A[4][56] ), .ip2(n12584), .op(n11973) );
  and2_1 U14932 ( .ip1(n12581), .ip2(\cache_data_A[7][56] ), .op(n11970) );
  nand2_1 U14933 ( .ip1(n12429), .ip2(\cache_data_A[6][56] ), .op(n11968) );
  nand2_1 U14934 ( .ip1(n12591), .ip2(\cache_data_A[3][56] ), .op(n11967) );
  nand2_1 U14935 ( .ip1(n12242), .ip2(\cache_data_A[1][56] ), .op(n11966) );
  nand2_1 U14936 ( .ip1(n11142), .ip2(\cache_data_A[2][56] ), .op(n11965) );
  nand4_1 U14937 ( .ip1(n11968), .ip2(n11967), .ip3(n11966), .ip4(n11965), 
        .op(n11969) );
  not_ab_or_c_or_d U14938 ( .ip1(\cache_data_A[0][56] ), .ip2(n12297), .ip3(
        n11970), .ip4(n11969), .op(n11972) );
  nand2_1 U14939 ( .ip1(n12118), .ip2(\cache_data_A[5][56] ), .op(n11971) );
  nand3_1 U14940 ( .ip1(n11973), .ip2(n11972), .ip3(n11971), .op(n13047) );
  nand2_1 U14941 ( .ip1(n12595), .ip2(n13047), .op(n11974) );
  nand3_1 U14942 ( .ip1(n11976), .ip2(n11975), .ip3(n11974), .op(n11977) );
  mux2_1 U14943 ( .ip1(N4132), .ip2(n11977), .s(n12599), .op(n5296) );
  nand2_1 U14944 ( .ip1(n12591), .ip2(\cache_data_A[3][121] ), .op(n11986) );
  and2_1 U14945 ( .ip1(n12581), .ip2(\cache_data_A[7][121] ), .op(n11983) );
  nand2_1 U14946 ( .ip1(n12429), .ip2(\cache_data_A[6][121] ), .op(n11981) );
  nand2_1 U14947 ( .ip1(n12475), .ip2(\cache_data_A[2][121] ), .op(n11980) );
  nand2_1 U14948 ( .ip1(n12582), .ip2(\cache_data_A[5][121] ), .op(n11979) );
  nand2_1 U14949 ( .ip1(n12476), .ip2(\cache_data_A[4][121] ), .op(n11978) );
  nand4_1 U14950 ( .ip1(n11981), .ip2(n11980), .ip3(n11979), .ip4(n11978), 
        .op(n11982) );
  not_ab_or_c_or_d U14951 ( .ip1(\cache_data_A[0][121] ), .ip2(n12297), .ip3(
        n11983), .ip4(n11982), .op(n11985) );
  nand2_1 U14952 ( .ip1(n12242), .ip2(\cache_data_A[1][121] ), .op(n11984) );
  nand3_1 U14953 ( .ip1(n11986), .ip2(n11985), .ip3(n11984), .op(n13065) );
  nand2_1 U14954 ( .ip1(n12509), .ip2(n13065), .op(n12060) );
  nand2_1 U14955 ( .ip1(n11057), .ip2(\cache_data_B[7][121] ), .op(n11995) );
  and2_1 U14956 ( .ip1(n11724), .ip2(\cache_data_B[1][121] ), .op(n11992) );
  nand2_1 U14957 ( .ip1(n11855), .ip2(\cache_data_B[2][121] ), .op(n11990) );
  nand2_1 U14958 ( .ip1(n12429), .ip2(\cache_data_B[6][121] ), .op(n11989) );
  nand2_1 U14959 ( .ip1(n12582), .ip2(\cache_data_B[5][121] ), .op(n11988) );
  nand2_1 U14960 ( .ip1(n12297), .ip2(\cache_data_B[0][121] ), .op(n11987) );
  nand4_1 U14961 ( .ip1(n11990), .ip2(n11989), .ip3(n11988), .ip4(n11987), 
        .op(n11991) );
  not_ab_or_c_or_d U14962 ( .ip1(n12096), .ip2(\cache_data_B[3][121] ), .ip3(
        n11992), .ip4(n11991), .op(n11994) );
  nand2_1 U14963 ( .ip1(n12194), .ip2(\cache_data_B[4][121] ), .op(n11993) );
  nand3_1 U14964 ( .ip1(n11995), .ip2(n11994), .ip3(n11993), .op(n13066) );
  nand2_1 U14965 ( .ip1(n12475), .ip2(\cache_data_A[2][89] ), .op(n11999) );
  nand2_1 U14966 ( .ip1(n10702), .ip2(\cache_data_A[7][89] ), .op(n11998) );
  nand2_1 U14967 ( .ip1(n12242), .ip2(\cache_data_A[1][89] ), .op(n11997) );
  nand2_1 U14968 ( .ip1(n12429), .ip2(\cache_data_A[6][89] ), .op(n11996) );
  nand4_1 U14969 ( .ip1(n11999), .ip2(n11998), .ip3(n11997), .ip4(n11996), 
        .op(n12005) );
  nand2_1 U14970 ( .ip1(n12297), .ip2(\cache_data_A[0][89] ), .op(n12003) );
  nand2_1 U14971 ( .ip1(n12194), .ip2(\cache_data_A[4][89] ), .op(n12002) );
  nand2_1 U14972 ( .ip1(n12591), .ip2(\cache_data_A[3][89] ), .op(n12001) );
  nand2_1 U14973 ( .ip1(n12582), .ip2(\cache_data_A[5][89] ), .op(n12000) );
  nand4_1 U14974 ( .ip1(n12003), .ip2(n12002), .ip3(n12001), .ip4(n12000), 
        .op(n12004) );
  nor2_1 U14975 ( .ip1(n12005), .ip2(n12004), .op(n13054) );
  nor2_1 U14976 ( .ip1(n13054), .ip2(n12529), .op(n12047) );
  nand2_1 U14977 ( .ip1(\cache_data_A[7][25] ), .ip2(n12552), .op(n12014) );
  and2_1 U14978 ( .ip1(n12591), .ip2(\cache_data_A[3][25] ), .op(n12011) );
  nand2_1 U14979 ( .ip1(n12475), .ip2(\cache_data_A[2][25] ), .op(n12009) );
  nand2_1 U14980 ( .ip1(n12582), .ip2(\cache_data_A[5][25] ), .op(n12008) );
  nand2_1 U14981 ( .ip1(n11156), .ip2(\cache_data_A[4][25] ), .op(n12007) );
  nand2_1 U14982 ( .ip1(n12204), .ip2(\cache_data_A[0][25] ), .op(n12006) );
  nand4_1 U14983 ( .ip1(n12009), .ip2(n12008), .ip3(n12007), .ip4(n12006), 
        .op(n12010) );
  not_ab_or_c_or_d U14984 ( .ip1(\cache_data_A[6][25] ), .ip2(n12337), .ip3(
        n12011), .ip4(n12010), .op(n12013) );
  nand2_1 U14985 ( .ip1(n12242), .ip2(\cache_data_A[1][25] ), .op(n12012) );
  nand3_1 U14986 ( .ip1(n12014), .ip2(n12013), .ip3(n12012), .op(n13056) );
  nand2_1 U14987 ( .ip1(n12550), .ip2(n13056), .op(n12045) );
  nand2_1 U14988 ( .ip1(\cache_data_B[0][57] ), .ip2(n12204), .op(n12023) );
  and2_1 U14989 ( .ip1(n12396), .ip2(\cache_data_B[4][57] ), .op(n12020) );
  nand2_1 U14990 ( .ip1(n10702), .ip2(\cache_data_B[7][57] ), .op(n12018) );
  nand2_1 U14991 ( .ip1(n12591), .ip2(\cache_data_B[3][57] ), .op(n12017) );
  nand2_1 U14992 ( .ip1(n12475), .ip2(\cache_data_B[2][57] ), .op(n12016) );
  nand2_1 U14993 ( .ip1(n12256), .ip2(\cache_data_B[5][57] ), .op(n12015) );
  nand4_1 U14994 ( .ip1(n12018), .ip2(n12017), .ip3(n12016), .ip4(n12015), 
        .op(n12019) );
  not_ab_or_c_or_d U14995 ( .ip1(\cache_data_B[6][57] ), .ip2(n12551), .ip3(
        n12020), .ip4(n12019), .op(n12022) );
  nand2_1 U14996 ( .ip1(n12242), .ip2(\cache_data_B[1][57] ), .op(n12021) );
  nand3_1 U14997 ( .ip1(n12023), .ip2(n12022), .ip3(n12021), .op(n13053) );
  nand2_1 U14998 ( .ip1(n12563), .ip2(n13053), .op(n12044) );
  nand2_1 U14999 ( .ip1(n12475), .ip2(\cache_data_B[2][25] ), .op(n12032) );
  and2_1 U15000 ( .ip1(n12468), .ip2(\cache_data_B[7][25] ), .op(n12029) );
  nand2_1 U15001 ( .ip1(n12582), .ip2(\cache_data_B[5][25] ), .op(n12027) );
  nand2_1 U15002 ( .ip1(n12242), .ip2(\cache_data_B[1][25] ), .op(n12026) );
  nand2_1 U15003 ( .ip1(n12591), .ip2(\cache_data_B[3][25] ), .op(n12025) );
  nand2_1 U15004 ( .ip1(n12429), .ip2(\cache_data_B[6][25] ), .op(n12024) );
  nand4_1 U15005 ( .ip1(n12027), .ip2(n12026), .ip3(n12025), .ip4(n12024), 
        .op(n12028) );
  not_ab_or_c_or_d U15006 ( .ip1(\cache_data_B[0][25] ), .ip2(n12297), .ip3(
        n12029), .ip4(n12028), .op(n12031) );
  nand2_1 U15007 ( .ip1(n11156), .ip2(\cache_data_B[4][25] ), .op(n12030) );
  nand3_1 U15008 ( .ip1(n12032), .ip2(n12031), .ip3(n12030), .op(n13055) );
  nand2_1 U15009 ( .ip1(n12539), .ip2(n13055), .op(n12043) );
  nand2_1 U15010 ( .ip1(n12476), .ip2(\cache_data_A[4][57] ), .op(n12041) );
  and2_1 U15011 ( .ip1(n12591), .ip2(\cache_data_A[3][57] ), .op(n12038) );
  nand2_1 U15012 ( .ip1(n12242), .ip2(\cache_data_A[1][57] ), .op(n12036) );
  nand2_1 U15013 ( .ip1(n12429), .ip2(\cache_data_A[6][57] ), .op(n12035) );
  nand2_1 U15014 ( .ip1(n12204), .ip2(\cache_data_A[0][57] ), .op(n12034) );
  nand2_1 U15015 ( .ip1(n11057), .ip2(\cache_data_A[7][57] ), .op(n12033) );
  nand4_1 U15016 ( .ip1(n12036), .ip2(n12035), .ip3(n12034), .ip4(n12033), 
        .op(n12037) );
  not_ab_or_c_or_d U15017 ( .ip1(\cache_data_A[2][57] ), .ip2(n12546), .ip3(
        n12038), .ip4(n12037), .op(n12040) );
  nand2_1 U15018 ( .ip1(n12582), .ip2(\cache_data_A[5][57] ), .op(n12039) );
  nand3_1 U15019 ( .ip1(n12041), .ip2(n12040), .ip3(n12039), .op(n13057) );
  nand2_1 U15020 ( .ip1(n12595), .ip2(n13057), .op(n12042) );
  nand4_1 U15021 ( .ip1(n12045), .ip2(n12044), .ip3(n12043), .ip4(n12042), 
        .op(n12046) );
  not_ab_or_c_or_d U15022 ( .ip1(n12573), .ip2(n13066), .ip3(n12047), .ip4(
        n12046), .op(n12059) );
  nand2_1 U15023 ( .ip1(n12475), .ip2(\cache_data_B[2][89] ), .op(n12057) );
  and2_1 U15024 ( .ip1(n12147), .ip2(\cache_data_B[1][89] ), .op(n12053) );
  nand2_1 U15025 ( .ip1(n8452), .ip2(\cache_data_B[0][89] ), .op(n12051) );
  nand2_1 U15026 ( .ip1(n12582), .ip2(\cache_data_B[5][89] ), .op(n12050) );
  nand2_1 U15027 ( .ip1(n12551), .ip2(\cache_data_B[6][89] ), .op(n12049) );
  nand2_1 U15028 ( .ip1(n10702), .ip2(\cache_data_B[7][89] ), .op(n12048) );
  nand4_1 U15029 ( .ip1(n12051), .ip2(n12050), .ip3(n12049), .ip4(n12048), 
        .op(n12052) );
  not_ab_or_c_or_d U15030 ( .ip1(\cache_data_B[4][89] ), .ip2(n12054), .ip3(
        n12053), .ip4(n12052), .op(n12056) );
  nand2_1 U15031 ( .ip1(n12591), .ip2(\cache_data_B[3][89] ), .op(n12055) );
  nand3_1 U15032 ( .ip1(n12057), .ip2(n12056), .ip3(n12055), .op(n13058) );
  nand2_1 U15033 ( .ip1(n12580), .ip2(n13058), .op(n12058) );
  nand3_1 U15034 ( .ip1(n12060), .ip2(n12059), .ip3(n12058), .op(n12061) );
  mux2_1 U15035 ( .ip1(N4129), .ip2(n12061), .s(n12599), .op(n5295) );
  nand2_1 U15036 ( .ip1(n12357), .ip2(\cache_data_B[0][90] ), .op(n12070) );
  and2_1 U15037 ( .ip1(n12468), .ip2(\cache_data_B[7][90] ), .op(n12067) );
  nand2_1 U15038 ( .ip1(n12242), .ip2(\cache_data_B[1][90] ), .op(n12065) );
  nand2_1 U15039 ( .ip1(n12591), .ip2(\cache_data_B[3][90] ), .op(n12064) );
  nand2_1 U15040 ( .ip1(n11156), .ip2(\cache_data_B[4][90] ), .op(n12063) );
  nand2_1 U15041 ( .ip1(n12582), .ip2(\cache_data_B[5][90] ), .op(n12062) );
  nand4_1 U15042 ( .ip1(n12065), .ip2(n12064), .ip3(n12063), .ip4(n12062), 
        .op(n12066) );
  not_ab_or_c_or_d U15043 ( .ip1(\cache_data_B[2][90] ), .ip2(n12546), .ip3(
        n12067), .ip4(n12066), .op(n12069) );
  nand2_1 U15044 ( .ip1(n12320), .ip2(\cache_data_B[6][90] ), .op(n12068) );
  nand3_1 U15045 ( .ip1(n12070), .ip2(n12069), .ip3(n12068), .op(n13071) );
  nand2_1 U15046 ( .ip1(n12580), .ip2(n13071), .op(n12145) );
  nand2_1 U15047 ( .ip1(n12475), .ip2(\cache_data_A[2][26] ), .op(n12079) );
  and2_1 U15048 ( .ip1(n12147), .ip2(\cache_data_A[1][26] ), .op(n12076) );
  nand2_1 U15049 ( .ip1(n12118), .ip2(\cache_data_A[5][26] ), .op(n12074) );
  nand2_1 U15050 ( .ip1(n10575), .ip2(\cache_data_A[7][26] ), .op(n12073) );
  nand2_1 U15051 ( .ip1(n12591), .ip2(\cache_data_A[3][26] ), .op(n12072) );
  nand2_1 U15052 ( .ip1(n11156), .ip2(\cache_data_A[4][26] ), .op(n12071) );
  nand4_1 U15053 ( .ip1(n12074), .ip2(n12073), .ip3(n12072), .ip4(n12071), 
        .op(n12075) );
  not_ab_or_c_or_d U15054 ( .ip1(n8452), .ip2(\cache_data_A[0][26] ), .ip3(
        n12076), .ip4(n12075), .op(n12078) );
  nand2_1 U15055 ( .ip1(n12320), .ip2(\cache_data_A[6][26] ), .op(n12077) );
  nand3_1 U15056 ( .ip1(n12079), .ip2(n12078), .ip3(n12077), .op(n13075) );
  nand2_1 U15057 ( .ip1(n12552), .ip2(\cache_data_A[7][90] ), .op(n12083) );
  nand2_1 U15058 ( .ip1(n8452), .ip2(\cache_data_A[0][90] ), .op(n12082) );
  nand2_1 U15059 ( .ip1(n12320), .ip2(\cache_data_A[6][90] ), .op(n12081) );
  nand2_1 U15060 ( .ip1(n12475), .ip2(\cache_data_A[2][90] ), .op(n12080) );
  nand4_1 U15061 ( .ip1(n12083), .ip2(n12082), .ip3(n12081), .ip4(n12080), 
        .op(n12089) );
  nand2_1 U15062 ( .ip1(n12256), .ip2(\cache_data_A[5][90] ), .op(n12087) );
  nand2_1 U15063 ( .ip1(n12242), .ip2(\cache_data_A[1][90] ), .op(n12086) );
  nand2_1 U15064 ( .ip1(n12591), .ip2(\cache_data_A[3][90] ), .op(n12085) );
  nand2_1 U15065 ( .ip1(n12396), .ip2(\cache_data_A[4][90] ), .op(n12084) );
  nand4_1 U15066 ( .ip1(n12087), .ip2(n12086), .ip3(n12085), .ip4(n12084), 
        .op(n12088) );
  nor2_1 U15067 ( .ip1(n12089), .ip2(n12088), .op(n13072) );
  nor2_1 U15068 ( .ip1(n13072), .ip2(n12529), .op(n12133) );
  nand2_1 U15069 ( .ip1(\cache_data_B[0][122] ), .ip2(n12204), .op(n12099) );
  and2_1 U15070 ( .ip1(n11280), .ip2(\cache_data_B[5][122] ), .op(n12095) );
  nand2_1 U15071 ( .ip1(n10702), .ip2(\cache_data_B[7][122] ), .op(n12093) );
  nand2_1 U15072 ( .ip1(n12320), .ip2(\cache_data_B[6][122] ), .op(n12092) );
  nand2_1 U15073 ( .ip1(n12396), .ip2(\cache_data_B[4][122] ), .op(n12091) );
  nand2_1 U15074 ( .ip1(n12242), .ip2(\cache_data_B[1][122] ), .op(n12090) );
  nand4_1 U15075 ( .ip1(n12093), .ip2(n12092), .ip3(n12091), .ip4(n12090), 
        .op(n12094) );
  not_ab_or_c_or_d U15076 ( .ip1(n12096), .ip2(\cache_data_B[3][122] ), .ip3(
        n12095), .ip4(n12094), .op(n12098) );
  nand2_1 U15077 ( .ip1(n11142), .ip2(\cache_data_B[2][122] ), .op(n12097) );
  nand3_1 U15078 ( .ip1(n12099), .ip2(n12098), .ip3(n12097), .op(n13076) );
  nand2_1 U15079 ( .ip1(n12573), .ip2(n13076), .op(n12131) );
  nand2_1 U15080 ( .ip1(n8452), .ip2(\cache_data_B[0][26] ), .op(n12108) );
  and2_1 U15081 ( .ip1(n12256), .ip2(\cache_data_B[5][26] ), .op(n12105) );
  nand2_1 U15082 ( .ip1(n12242), .ip2(\cache_data_B[1][26] ), .op(n12103) );
  nand2_1 U15083 ( .ip1(n11057), .ip2(\cache_data_B[7][26] ), .op(n12102) );
  nand2_1 U15084 ( .ip1(n12396), .ip2(\cache_data_B[4][26] ), .op(n12101) );
  nand2_1 U15085 ( .ip1(n12475), .ip2(\cache_data_B[2][26] ), .op(n12100) );
  nand4_1 U15086 ( .ip1(n12103), .ip2(n12102), .ip3(n12101), .ip4(n12100), 
        .op(n12104) );
  not_ab_or_c_or_d U15087 ( .ip1(\cache_data_B[3][26] ), .ip2(n12559), .ip3(
        n12105), .ip4(n12104), .op(n12107) );
  nand2_1 U15088 ( .ip1(n12320), .ip2(\cache_data_B[6][26] ), .op(n12106) );
  nand3_1 U15089 ( .ip1(n12108), .ip2(n12107), .ip3(n12106), .op(n13083) );
  nand2_1 U15090 ( .ip1(n12539), .ip2(n13083), .op(n12130) );
  nand2_1 U15091 ( .ip1(n12552), .ip2(\cache_data_B[7][58] ), .op(n12117) );
  and2_1 U15092 ( .ip1(n11156), .ip2(\cache_data_B[4][58] ), .op(n12114) );
  nand2_1 U15093 ( .ip1(n12582), .ip2(\cache_data_B[5][58] ), .op(n12112) );
  nand2_1 U15094 ( .ip1(n12204), .ip2(\cache_data_B[0][58] ), .op(n12111) );
  nand2_1 U15095 ( .ip1(n12242), .ip2(\cache_data_B[1][58] ), .op(n12110) );
  nand2_1 U15096 ( .ip1(n12591), .ip2(\cache_data_B[3][58] ), .op(n12109) );
  nand4_1 U15097 ( .ip1(n12112), .ip2(n12111), .ip3(n12110), .ip4(n12109), 
        .op(n12113) );
  not_ab_or_c_or_d U15098 ( .ip1(n12546), .ip2(\cache_data_B[2][58] ), .ip3(
        n12114), .ip4(n12113), .op(n12116) );
  nand2_1 U15099 ( .ip1(n12320), .ip2(\cache_data_B[6][58] ), .op(n12115) );
  nand3_1 U15100 ( .ip1(n12117), .ip2(n12116), .ip3(n12115), .op(n13084) );
  nand2_1 U15101 ( .ip1(n12563), .ip2(n13084), .op(n12129) );
  nand2_1 U15102 ( .ip1(n10702), .ip2(\cache_data_A[7][122] ), .op(n12127) );
  and2_1 U15103 ( .ip1(n12486), .ip2(\cache_data_A[2][122] ), .op(n12124) );
  nand2_1 U15104 ( .ip1(n12118), .ip2(\cache_data_A[5][122] ), .op(n12122) );
  nand2_1 U15105 ( .ip1(n11324), .ip2(\cache_data_A[4][122] ), .op(n12121) );
  nand2_1 U15106 ( .ip1(n12320), .ip2(\cache_data_A[6][122] ), .op(n12120) );
  nand2_1 U15107 ( .ip1(n12591), .ip2(\cache_data_A[3][122] ), .op(n12119) );
  nand4_1 U15108 ( .ip1(n12122), .ip2(n12121), .ip3(n12120), .ip4(n12119), 
        .op(n12123) );
  not_ab_or_c_or_d U15109 ( .ip1(n11911), .ip2(\cache_data_A[0][122] ), .ip3(
        n12124), .ip4(n12123), .op(n12126) );
  nand2_1 U15110 ( .ip1(n12242), .ip2(\cache_data_A[1][122] ), .op(n12125) );
  nand3_1 U15111 ( .ip1(n12127), .ip2(n12126), .ip3(n12125), .op(n13074) );
  nand2_1 U15112 ( .ip1(n12509), .ip2(n13074), .op(n12128) );
  nand4_1 U15113 ( .ip1(n12131), .ip2(n12130), .ip3(n12129), .ip4(n12128), 
        .op(n12132) );
  not_ab_or_c_or_d U15114 ( .ip1(n12550), .ip2(n13075), .ip3(n12133), .ip4(
        n12132), .op(n12144) );
  nand2_1 U15115 ( .ip1(\cache_data_A[0][58] ), .ip2(n12370), .op(n12142) );
  and2_1 U15116 ( .ip1(n12429), .ip2(\cache_data_A[6][58] ), .op(n12139) );
  nand2_1 U15117 ( .ip1(n12591), .ip2(\cache_data_A[3][58] ), .op(n12137) );
  nand2_1 U15118 ( .ip1(n12582), .ip2(\cache_data_A[5][58] ), .op(n12136) );
  nand2_1 U15119 ( .ip1(n12396), .ip2(\cache_data_A[4][58] ), .op(n12135) );
  nand2_1 U15120 ( .ip1(n12242), .ip2(\cache_data_A[1][58] ), .op(n12134) );
  nand4_1 U15121 ( .ip1(n12137), .ip2(n12136), .ip3(n12135), .ip4(n12134), 
        .op(n12138) );
  not_ab_or_c_or_d U15122 ( .ip1(\cache_data_A[2][58] ), .ip2(n12546), .ip3(
        n12139), .ip4(n12138), .op(n12141) );
  nand2_1 U15123 ( .ip1(n10702), .ip2(\cache_data_A[7][58] ), .op(n12140) );
  nand3_1 U15124 ( .ip1(n12142), .ip2(n12141), .ip3(n12140), .op(n13073) );
  nand2_1 U15125 ( .ip1(n12595), .ip2(n13073), .op(n12143) );
  nand3_1 U15126 ( .ip1(n12145), .ip2(n12144), .ip3(n12143), .op(n12146) );
  mux2_1 U15127 ( .ip1(N4126), .ip2(n12146), .s(n12599), .op(n5294) );
  nand2_1 U15128 ( .ip1(\cache_data_A[0][123] ), .ip2(n12370), .op(n12156) );
  and2_1 U15129 ( .ip1(n12147), .ip2(\cache_data_A[1][123] ), .op(n12153) );
  nand2_1 U15130 ( .ip1(n12582), .ip2(\cache_data_A[5][123] ), .op(n12151) );
  nand2_1 U15131 ( .ip1(n12475), .ip2(\cache_data_A[2][123] ), .op(n12150) );
  nand2_1 U15132 ( .ip1(n11057), .ip2(\cache_data_A[7][123] ), .op(n12149) );
  nand2_1 U15133 ( .ip1(n12591), .ip2(\cache_data_A[3][123] ), .op(n12148) );
  nand4_1 U15134 ( .ip1(n12151), .ip2(n12150), .ip3(n12149), .ip4(n12148), 
        .op(n12152) );
  not_ab_or_c_or_d U15135 ( .ip1(\cache_data_A[4][123] ), .ip2(n11156), .ip3(
        n12153), .ip4(n12152), .op(n12155) );
  nand2_1 U15136 ( .ip1(n12320), .ip2(\cache_data_A[6][123] ), .op(n12154) );
  nand3_1 U15137 ( .ip1(n12156), .ip2(n12155), .ip3(n12154), .op(n13092) );
  nand2_1 U15138 ( .ip1(n12509), .ip2(n13092), .op(n12231) );
  nand2_1 U15139 ( .ip1(n12552), .ip2(\cache_data_B[7][27] ), .op(n12165) );
  and2_1 U15140 ( .ip1(n10686), .ip2(\cache_data_B[1][27] ), .op(n12162) );
  nand2_1 U15141 ( .ip1(n12297), .ip2(\cache_data_B[0][27] ), .op(n12160) );
  nand2_1 U15142 ( .ip1(n12321), .ip2(\cache_data_B[3][27] ), .op(n12159) );
  nand2_1 U15143 ( .ip1(n12320), .ip2(\cache_data_B[6][27] ), .op(n12158) );
  nand2_1 U15144 ( .ip1(n12256), .ip2(\cache_data_B[5][27] ), .op(n12157) );
  nand4_1 U15145 ( .ip1(n12160), .ip2(n12159), .ip3(n12158), .ip4(n12157), 
        .op(n12161) );
  not_ab_or_c_or_d U15146 ( .ip1(\cache_data_B[2][27] ), .ip2(n12546), .ip3(
        n12162), .ip4(n12161), .op(n12164) );
  nand2_1 U15147 ( .ip1(n12396), .ip2(\cache_data_B[4][27] ), .op(n12163) );
  nand3_1 U15148 ( .ip1(n12165), .ip2(n12164), .ip3(n12163), .op(n13094) );
  nand2_1 U15149 ( .ip1(n12320), .ip2(\cache_data_A[6][91] ), .op(n12169) );
  nand2_1 U15150 ( .ip1(n12581), .ip2(\cache_data_A[7][91] ), .op(n12168) );
  nand2_1 U15151 ( .ip1(n12256), .ip2(\cache_data_A[5][91] ), .op(n12167) );
  nand2_1 U15152 ( .ip1(n8452), .ip2(\cache_data_A[0][91] ), .op(n12166) );
  nand4_1 U15153 ( .ip1(n12169), .ip2(n12168), .ip3(n12167), .ip4(n12166), 
        .op(n12175) );
  nand2_1 U15154 ( .ip1(n12410), .ip2(\cache_data_A[3][91] ), .op(n12173) );
  nand2_1 U15155 ( .ip1(n12475), .ip2(\cache_data_A[2][91] ), .op(n12172) );
  nand2_1 U15156 ( .ip1(n12242), .ip2(\cache_data_A[1][91] ), .op(n12171) );
  nand2_1 U15157 ( .ip1(n12396), .ip2(\cache_data_A[4][91] ), .op(n12170) );
  nand4_1 U15158 ( .ip1(n12173), .ip2(n12172), .ip3(n12171), .ip4(n12170), 
        .op(n12174) );
  nor2_1 U15159 ( .ip1(n12175), .ip2(n12174), .op(n13090) );
  nor2_1 U15160 ( .ip1(n13090), .ip2(n12529), .op(n12219) );
  nand2_1 U15161 ( .ip1(n12410), .ip2(\cache_data_B[3][91] ), .op(n12184) );
  and2_1 U15162 ( .ip1(n12256), .ip2(\cache_data_B[5][91] ), .op(n12181) );
  nand2_1 U15163 ( .ip1(n11057), .ip2(\cache_data_B[7][91] ), .op(n12179) );
  nand2_1 U15164 ( .ip1(n12320), .ip2(\cache_data_B[6][91] ), .op(n12178) );
  nand2_1 U15165 ( .ip1(n8452), .ip2(\cache_data_B[0][91] ), .op(n12177) );
  nand2_1 U15166 ( .ip1(n12242), .ip2(\cache_data_B[1][91] ), .op(n12176) );
  nand4_1 U15167 ( .ip1(n12179), .ip2(n12178), .ip3(n12177), .ip4(n12176), 
        .op(n12180) );
  not_ab_or_c_or_d U15168 ( .ip1(\cache_data_B[2][91] ), .ip2(n12546), .ip3(
        n12181), .ip4(n12180), .op(n12183) );
  nand2_1 U15169 ( .ip1(n12396), .ip2(\cache_data_B[4][91] ), .op(n12182) );
  nand3_1 U15170 ( .ip1(n12184), .ip2(n12183), .ip3(n12182), .op(n13089) );
  nand2_1 U15171 ( .ip1(n12580), .ip2(n13089), .op(n12217) );
  nand2_1 U15172 ( .ip1(n12320), .ip2(\cache_data_B[6][59] ), .op(n12193) );
  and2_1 U15173 ( .ip1(n12256), .ip2(\cache_data_B[5][59] ), .op(n12190) );
  nand2_1 U15174 ( .ip1(n8452), .ip2(\cache_data_B[0][59] ), .op(n12188) );
  nand2_1 U15175 ( .ip1(n12475), .ip2(\cache_data_B[2][59] ), .op(n12187) );
  nand2_1 U15176 ( .ip1(n12396), .ip2(\cache_data_B[4][59] ), .op(n12186) );
  nand2_1 U15177 ( .ip1(n12410), .ip2(\cache_data_B[3][59] ), .op(n12185) );
  nand4_1 U15178 ( .ip1(n12188), .ip2(n12187), .ip3(n12186), .ip4(n12185), 
        .op(n12189) );
  not_ab_or_c_or_d U15179 ( .ip1(\cache_data_B[7][59] ), .ip2(n11057), .ip3(
        n12190), .ip4(n12189), .op(n12192) );
  nand2_1 U15180 ( .ip1(n12242), .ip2(\cache_data_B[1][59] ), .op(n12191) );
  nand3_1 U15181 ( .ip1(n12193), .ip2(n12192), .ip3(n12191), .op(n13101) );
  nand2_1 U15182 ( .ip1(n12563), .ip2(n13101), .op(n12216) );
  nand2_1 U15183 ( .ip1(n11855), .ip2(\cache_data_A[2][59] ), .op(n12203) );
  and2_1 U15184 ( .ip1(n12194), .ip2(\cache_data_A[4][59] ), .op(n12200) );
  nand2_1 U15185 ( .ip1(n12242), .ip2(\cache_data_A[1][59] ), .op(n12198) );
  nand2_1 U15186 ( .ip1(n11057), .ip2(\cache_data_A[7][59] ), .op(n12197) );
  nand2_1 U15187 ( .ip1(n12320), .ip2(\cache_data_A[6][59] ), .op(n12196) );
  nand2_1 U15188 ( .ip1(n12410), .ip2(\cache_data_A[3][59] ), .op(n12195) );
  nand4_1 U15189 ( .ip1(n12198), .ip2(n12197), .ip3(n12196), .ip4(n12195), 
        .op(n12199) );
  not_ab_or_c_or_d U15190 ( .ip1(\cache_data_A[0][59] ), .ip2(n12297), .ip3(
        n12200), .ip4(n12199), .op(n12202) );
  nand2_1 U15191 ( .ip1(n12256), .ip2(\cache_data_A[5][59] ), .op(n12201) );
  nand3_1 U15192 ( .ip1(n12203), .ip2(n12202), .ip3(n12201), .op(n13102) );
  nand2_1 U15193 ( .ip1(n12595), .ip2(n13102), .op(n12215) );
  nand2_1 U15194 ( .ip1(\cache_data_B[0][123] ), .ip2(n12204), .op(n12213) );
  and2_1 U15195 ( .ip1(n12371), .ip2(\cache_data_B[6][123] ), .op(n12210) );
  nand2_1 U15196 ( .ip1(n12410), .ip2(\cache_data_B[3][123] ), .op(n12208) );
  nand2_1 U15197 ( .ip1(n12256), .ip2(\cache_data_B[5][123] ), .op(n12207) );
  nand2_1 U15198 ( .ip1(n12242), .ip2(\cache_data_B[1][123] ), .op(n12206) );
  nand2_1 U15199 ( .ip1(n12475), .ip2(\cache_data_B[2][123] ), .op(n12205) );
  nand4_1 U15200 ( .ip1(n12208), .ip2(n12207), .ip3(n12206), .ip4(n12205), 
        .op(n12209) );
  not_ab_or_c_or_d U15201 ( .ip1(\cache_data_B[7][123] ), .ip2(n12468), .ip3(
        n12210), .ip4(n12209), .op(n12212) );
  nand2_1 U15202 ( .ip1(n12396), .ip2(\cache_data_B[4][123] ), .op(n12211) );
  nand3_1 U15203 ( .ip1(n12213), .ip2(n12212), .ip3(n12211), .op(n13091) );
  nand2_1 U15204 ( .ip1(n12573), .ip2(n13091), .op(n12214) );
  nand4_1 U15205 ( .ip1(n12217), .ip2(n12216), .ip3(n12215), .ip4(n12214), 
        .op(n12218) );
  not_ab_or_c_or_d U15206 ( .ip1(n12539), .ip2(n13094), .ip3(n12219), .ip4(
        n12218), .op(n12230) );
  nand2_1 U15207 ( .ip1(n12297), .ip2(\cache_data_A[0][27] ), .op(n12228) );
  and2_1 U15208 ( .ip1(n12396), .ip2(\cache_data_A[4][27] ), .op(n12225) );
  nand2_1 U15209 ( .ip1(n12321), .ip2(\cache_data_A[3][27] ), .op(n12223) );
  nand2_1 U15210 ( .ip1(n12475), .ip2(\cache_data_A[2][27] ), .op(n12222) );
  nand2_1 U15211 ( .ip1(n12320), .ip2(\cache_data_A[6][27] ), .op(n12221) );
  nand2_1 U15212 ( .ip1(n12242), .ip2(\cache_data_A[1][27] ), .op(n12220) );
  nand4_1 U15213 ( .ip1(n12223), .ip2(n12222), .ip3(n12221), .ip4(n12220), 
        .op(n12224) );
  not_ab_or_c_or_d U15214 ( .ip1(n12278), .ip2(\cache_data_A[7][27] ), .ip3(
        n12225), .ip4(n12224), .op(n12227) );
  nand2_1 U15215 ( .ip1(n12256), .ip2(\cache_data_A[5][27] ), .op(n12226) );
  nand3_1 U15216 ( .ip1(n12228), .ip2(n12227), .ip3(n12226), .op(n13093) );
  nand2_1 U15217 ( .ip1(n12550), .ip2(n13093), .op(n12229) );
  nand3_1 U15218 ( .ip1(n12231), .ip2(n12230), .ip3(n12229), .op(n12232) );
  mux2_1 U15219 ( .ip1(N4123), .ip2(n12232), .s(n12599), .op(n5293) );
  nand2_1 U15220 ( .ip1(n12429), .ip2(\cache_data_B[6][60] ), .op(n12241) );
  and2_1 U15221 ( .ip1(n8060), .ip2(\cache_data_B[3][60] ), .op(n12238) );
  nand2_1 U15222 ( .ip1(n12475), .ip2(\cache_data_B[2][60] ), .op(n12236) );
  nand2_1 U15223 ( .ip1(n12357), .ip2(\cache_data_B[0][60] ), .op(n12235) );
  nand2_1 U15224 ( .ip1(n12396), .ip2(\cache_data_B[4][60] ), .op(n12234) );
  nand2_1 U15225 ( .ip1(n12242), .ip2(\cache_data_B[1][60] ), .op(n12233) );
  nand4_1 U15226 ( .ip1(n12236), .ip2(n12235), .ip3(n12234), .ip4(n12233), 
        .op(n12237) );
  not_ab_or_c_or_d U15227 ( .ip1(\cache_data_B[7][60] ), .ip2(n10702), .ip3(
        n12238), .ip4(n12237), .op(n12240) );
  nand2_1 U15228 ( .ip1(n12256), .ip2(\cache_data_B[5][60] ), .op(n12239) );
  nand3_1 U15229 ( .ip1(n12241), .ip2(n12240), .ip3(n12239), .op(n13120) );
  nand2_1 U15230 ( .ip1(n12563), .ip2(n13120), .op(n12318) );
  nand2_1 U15231 ( .ip1(n12396), .ip2(\cache_data_A[4][124] ), .op(n12251) );
  and2_1 U15232 ( .ip1(n12486), .ip2(\cache_data_A[2][124] ), .op(n12248) );
  nand2_1 U15233 ( .ip1(n12242), .ip2(\cache_data_A[1][124] ), .op(n12246) );
  nand2_1 U15234 ( .ip1(n11057), .ip2(\cache_data_A[7][124] ), .op(n12245) );
  nand2_1 U15235 ( .ip1(n12429), .ip2(\cache_data_A[6][124] ), .op(n12244) );
  nand2_1 U15236 ( .ip1(n12410), .ip2(\cache_data_A[3][124] ), .op(n12243) );
  nand4_1 U15237 ( .ip1(n12246), .ip2(n12245), .ip3(n12244), .ip4(n12243), 
        .op(n12247) );
  not_ab_or_c_or_d U15238 ( .ip1(n12297), .ip2(\cache_data_A[0][124] ), .ip3(
        n12248), .ip4(n12247), .op(n12250) );
  nand2_1 U15239 ( .ip1(n12256), .ip2(\cache_data_A[5][124] ), .op(n12249) );
  nand3_1 U15240 ( .ip1(n12251), .ip2(n12250), .ip3(n12249), .op(n13110) );
  nand2_1 U15241 ( .ip1(n12429), .ip2(\cache_data_A[6][92] ), .op(n12255) );
  nand2_1 U15242 ( .ip1(n12396), .ip2(\cache_data_A[4][92] ), .op(n12254) );
  nand2_1 U15243 ( .ip1(n12321), .ip2(\cache_data_A[3][92] ), .op(n12253) );
  nand2_1 U15244 ( .ip1(n12475), .ip2(\cache_data_A[2][92] ), .op(n12252) );
  nand4_1 U15245 ( .ip1(n12255), .ip2(n12254), .ip3(n12253), .ip4(n12252), 
        .op(n12262) );
  nand2_1 U15246 ( .ip1(n12581), .ip2(\cache_data_A[7][92] ), .op(n12260) );
  nand2_1 U15247 ( .ip1(n11946), .ip2(\cache_data_A[1][92] ), .op(n12259) );
  nand2_1 U15248 ( .ip1(n12297), .ip2(\cache_data_A[0][92] ), .op(n12258) );
  nand2_1 U15249 ( .ip1(n12256), .ip2(\cache_data_A[5][92] ), .op(n12257) );
  nand4_1 U15250 ( .ip1(n12260), .ip2(n12259), .ip3(n12258), .ip4(n12257), 
        .op(n12261) );
  nor2_1 U15251 ( .ip1(n12262), .ip2(n12261), .op(n13108) );
  nor2_1 U15252 ( .ip1(n13108), .ip2(n12529), .op(n12306) );
  nand2_1 U15253 ( .ip1(n8452), .ip2(\cache_data_B[0][124] ), .op(n12271) );
  and2_1 U15254 ( .ip1(n12396), .ip2(\cache_data_B[4][124] ), .op(n12268) );
  nand2_1 U15255 ( .ip1(n12458), .ip2(\cache_data_B[6][124] ), .op(n12266) );
  nand2_1 U15256 ( .ip1(n12475), .ip2(\cache_data_B[2][124] ), .op(n12265) );
  nand2_1 U15257 ( .ip1(n11280), .ip2(\cache_data_B[5][124] ), .op(n12264) );
  nand2_1 U15258 ( .ip1(n12410), .ip2(\cache_data_B[3][124] ), .op(n12263) );
  nand4_1 U15259 ( .ip1(n12266), .ip2(n12265), .ip3(n12264), .ip4(n12263), 
        .op(n12267) );
  not_ab_or_c_or_d U15260 ( .ip1(n12278), .ip2(\cache_data_B[7][124] ), .ip3(
        n12268), .ip4(n12267), .op(n12270) );
  nand2_1 U15261 ( .ip1(n11311), .ip2(\cache_data_B[1][124] ), .op(n12269) );
  nand3_1 U15262 ( .ip1(n12271), .ip2(n12270), .ip3(n12269), .op(n13109) );
  nand2_1 U15263 ( .ip1(n12573), .ip2(n13109), .op(n12304) );
  nand2_1 U15264 ( .ip1(n12429), .ip2(\cache_data_A[6][28] ), .op(n12281) );
  and2_1 U15265 ( .ip1(n8060), .ip2(\cache_data_A[3][28] ), .op(n12277) );
  nand2_1 U15266 ( .ip1(n8452), .ip2(\cache_data_A[0][28] ), .op(n12275) );
  nand2_1 U15267 ( .ip1(n12475), .ip2(\cache_data_A[2][28] ), .op(n12274) );
  nand2_1 U15268 ( .ip1(n12054), .ip2(\cache_data_A[4][28] ), .op(n12273) );
  nand2_1 U15269 ( .ip1(n11304), .ip2(\cache_data_A[5][28] ), .op(n12272) );
  nand4_1 U15270 ( .ip1(n12275), .ip2(n12274), .ip3(n12273), .ip4(n12272), 
        .op(n12276) );
  not_ab_or_c_or_d U15271 ( .ip1(\cache_data_A[7][28] ), .ip2(n12278), .ip3(
        n12277), .ip4(n12276), .op(n12280) );
  nand2_1 U15272 ( .ip1(n11946), .ip2(\cache_data_A[1][28] ), .op(n12279) );
  nand3_1 U15273 ( .ip1(n12281), .ip2(n12280), .ip3(n12279), .op(n13111) );
  nand2_1 U15274 ( .ip1(n12550), .ip2(n13111), .op(n12303) );
  nand2_1 U15275 ( .ip1(n12297), .ip2(\cache_data_B[0][92] ), .op(n12290) );
  and2_1 U15276 ( .ip1(n10686), .ip2(\cache_data_B[1][92] ), .op(n12287) );
  nand2_1 U15277 ( .ip1(n12410), .ip2(\cache_data_B[3][92] ), .op(n12285) );
  nand2_1 U15278 ( .ip1(n12475), .ip2(\cache_data_B[2][92] ), .op(n12284) );
  nand2_1 U15279 ( .ip1(n12396), .ip2(\cache_data_B[4][92] ), .op(n12283) );
  nand2_1 U15280 ( .ip1(n11304), .ip2(\cache_data_B[5][92] ), .op(n12282) );
  nand4_1 U15281 ( .ip1(n12285), .ip2(n12284), .ip3(n12283), .ip4(n12282), 
        .op(n12286) );
  not_ab_or_c_or_d U15282 ( .ip1(\cache_data_B[6][92] ), .ip2(n12337), .ip3(
        n12287), .ip4(n12286), .op(n12289) );
  nand2_1 U15283 ( .ip1(n12552), .ip2(\cache_data_B[7][92] ), .op(n12288) );
  nand3_1 U15284 ( .ip1(n12290), .ip2(n12289), .ip3(n12288), .op(n13107) );
  nand2_1 U15285 ( .ip1(n12580), .ip2(n13107), .op(n12302) );
  nand2_1 U15286 ( .ip1(\cache_data_A[2][60] ), .ip2(n12486), .op(n12300) );
  and2_1 U15287 ( .ip1(n12591), .ip2(\cache_data_A[3][60] ), .op(n12296) );
  nand2_1 U15288 ( .ip1(n12581), .ip2(\cache_data_A[7][60] ), .op(n12294) );
  nand2_1 U15289 ( .ip1(n12429), .ip2(\cache_data_A[6][60] ), .op(n12293) );
  nand2_1 U15290 ( .ip1(n12396), .ip2(\cache_data_A[4][60] ), .op(n12292) );
  nand2_1 U15291 ( .ip1(n11304), .ip2(\cache_data_A[5][60] ), .op(n12291) );
  nand4_1 U15292 ( .ip1(n12294), .ip2(n12293), .ip3(n12292), .ip4(n12291), 
        .op(n12295) );
  not_ab_or_c_or_d U15293 ( .ip1(n12297), .ip2(\cache_data_A[0][60] ), .ip3(
        n12296), .ip4(n12295), .op(n12299) );
  nand2_1 U15294 ( .ip1(n11946), .ip2(\cache_data_A[1][60] ), .op(n12298) );
  nand3_1 U15295 ( .ip1(n12300), .ip2(n12299), .ip3(n12298), .op(n13119) );
  nand2_1 U15296 ( .ip1(n12595), .ip2(n13119), .op(n12301) );
  nand4_1 U15297 ( .ip1(n12304), .ip2(n12303), .ip3(n12302), .ip4(n12301), 
        .op(n12305) );
  not_ab_or_c_or_d U15298 ( .ip1(n12509), .ip2(n13110), .ip3(n12306), .ip4(
        n12305), .op(n12317) );
  nand2_1 U15299 ( .ip1(n8452), .ip2(\cache_data_B[0][28] ), .op(n12315) );
  and2_1 U15300 ( .ip1(n12396), .ip2(\cache_data_B[4][28] ), .op(n12312) );
  nand2_1 U15301 ( .ip1(n12321), .ip2(\cache_data_B[3][28] ), .op(n12310) );
  nand2_1 U15302 ( .ip1(n11057), .ip2(\cache_data_B[7][28] ), .op(n12309) );
  nand2_1 U15303 ( .ip1(n10686), .ip2(\cache_data_B[1][28] ), .op(n12308) );
  nand2_1 U15304 ( .ip1(n11296), .ip2(\cache_data_B[5][28] ), .op(n12307) );
  nand4_1 U15305 ( .ip1(n12310), .ip2(n12309), .ip3(n12308), .ip4(n12307), 
        .op(n12311) );
  not_ab_or_c_or_d U15306 ( .ip1(n12551), .ip2(\cache_data_B[6][28] ), .ip3(
        n12312), .ip4(n12311), .op(n12314) );
  nand2_1 U15307 ( .ip1(n11855), .ip2(\cache_data_B[2][28] ), .op(n12313) );
  nand3_1 U15308 ( .ip1(n12315), .ip2(n12314), .ip3(n12313), .op(n13112) );
  nand2_1 U15309 ( .ip1(n12539), .ip2(n13112), .op(n12316) );
  nand3_1 U15310 ( .ip1(n12318), .ip2(n12317), .ip3(n12316), .op(n12319) );
  mux2_1 U15311 ( .ip1(N4120), .ip2(n12319), .s(n12599), .op(n5292) );
  nand2_1 U15312 ( .ip1(n10575), .ip2(\cache_data_B[7][125] ), .op(n12330) );
  and2_1 U15313 ( .ip1(n12147), .ip2(\cache_data_B[1][125] ), .op(n12327) );
  nand2_1 U15314 ( .ip1(n12475), .ip2(\cache_data_B[2][125] ), .op(n12325) );
  nand2_1 U15315 ( .ip1(n12320), .ip2(\cache_data_B[6][125] ), .op(n12324) );
  nand2_1 U15316 ( .ip1(n12297), .ip2(\cache_data_B[0][125] ), .op(n12323) );
  nand2_1 U15317 ( .ip1(n12321), .ip2(\cache_data_B[3][125] ), .op(n12322) );
  nand4_1 U15318 ( .ip1(n12325), .ip2(n12324), .ip3(n12323), .ip4(n12322), 
        .op(n12326) );
  not_ab_or_c_or_d U15319 ( .ip1(n12194), .ip2(\cache_data_B[4][125] ), .ip3(
        n12327), .ip4(n12326), .op(n12329) );
  nand2_1 U15320 ( .ip1(n12582), .ip2(\cache_data_B[5][125] ), .op(n12328) );
  nand3_1 U15321 ( .ip1(n12330), .ip2(n12329), .ip3(n12328), .op(n13125) );
  nand2_1 U15322 ( .ip1(n12573), .ip2(n13125), .op(n12408) );
  nand2_1 U15323 ( .ip1(\cache_data_A[0][125] ), .ip2(n12370), .op(n12340) );
  and2_1 U15324 ( .ip1(n12591), .ip2(\cache_data_A[3][125] ), .op(n12336) );
  nand2_1 U15325 ( .ip1(n12581), .ip2(\cache_data_A[7][125] ), .op(n12334) );
  nand2_1 U15326 ( .ip1(n12475), .ip2(\cache_data_A[2][125] ), .op(n12333) );
  nand2_1 U15327 ( .ip1(n12242), .ip2(\cache_data_A[1][125] ), .op(n12332) );
  nand2_1 U15328 ( .ip1(n11304), .ip2(\cache_data_A[5][125] ), .op(n12331) );
  nand4_1 U15329 ( .ip1(n12334), .ip2(n12333), .ip3(n12332), .ip4(n12331), 
        .op(n12335) );
  not_ab_or_c_or_d U15330 ( .ip1(\cache_data_A[6][125] ), .ip2(n12337), .ip3(
        n12336), .ip4(n12335), .op(n12339) );
  nand2_1 U15331 ( .ip1(n12476), .ip2(\cache_data_A[4][125] ), .op(n12338) );
  nand3_1 U15332 ( .ip1(n12340), .ip2(n12339), .ip3(n12338), .op(n13130) );
  nand2_1 U15333 ( .ip1(n8452), .ip2(\cache_data_A[0][93] ), .op(n12344) );
  nand2_1 U15334 ( .ip1(n12429), .ip2(\cache_data_A[6][93] ), .op(n12343) );
  nand2_1 U15335 ( .ip1(n12582), .ip2(\cache_data_A[5][93] ), .op(n12342) );
  nand2_1 U15336 ( .ip1(n12581), .ip2(\cache_data_A[7][93] ), .op(n12341) );
  nand4_1 U15337 ( .ip1(n12344), .ip2(n12343), .ip3(n12342), .ip4(n12341), 
        .op(n12350) );
  nand2_1 U15338 ( .ip1(n10686), .ip2(\cache_data_A[1][93] ), .op(n12348) );
  nand2_1 U15339 ( .ip1(n12476), .ip2(\cache_data_A[4][93] ), .op(n12347) );
  nand2_1 U15340 ( .ip1(n12475), .ip2(\cache_data_A[2][93] ), .op(n12346) );
  nand2_1 U15341 ( .ip1(n12410), .ip2(\cache_data_A[3][93] ), .op(n12345) );
  nand4_1 U15342 ( .ip1(n12348), .ip2(n12347), .ip3(n12346), .ip4(n12345), 
        .op(n12349) );
  nor2_1 U15343 ( .ip1(n12350), .ip2(n12349), .op(n13126) );
  nor2_1 U15344 ( .ip1(n13126), .ip2(n12529), .op(n12395) );
  nand2_1 U15345 ( .ip1(n12321), .ip2(\cache_data_B[3][29] ), .op(n12360) );
  and2_1 U15346 ( .ip1(n12486), .ip2(\cache_data_B[2][29] ), .op(n12356) );
  nand2_1 U15347 ( .ip1(n12429), .ip2(\cache_data_B[6][29] ), .op(n12354) );
  nand2_1 U15348 ( .ip1(n11057), .ip2(\cache_data_B[7][29] ), .op(n12353) );
  nand2_1 U15349 ( .ip1(n12242), .ip2(\cache_data_B[1][29] ), .op(n12352) );
  nand2_1 U15350 ( .ip1(n11280), .ip2(\cache_data_B[5][29] ), .op(n12351) );
  nand4_1 U15351 ( .ip1(n12354), .ip2(n12353), .ip3(n12352), .ip4(n12351), 
        .op(n12355) );
  not_ab_or_c_or_d U15352 ( .ip1(\cache_data_B[0][29] ), .ip2(n12357), .ip3(
        n12356), .ip4(n12355), .op(n12359) );
  nand2_1 U15353 ( .ip1(n12476), .ip2(\cache_data_B[4][29] ), .op(n12358) );
  nand3_1 U15354 ( .ip1(n12360), .ip2(n12359), .ip3(n12358), .op(n13127) );
  nand2_1 U15355 ( .ip1(n12539), .ip2(n13127), .op(n12393) );
  nand2_1 U15356 ( .ip1(n12476), .ip2(\cache_data_A[4][29] ), .op(n12369) );
  and2_1 U15357 ( .ip1(n12429), .ip2(\cache_data_A[6][29] ), .op(n12366) );
  nand2_1 U15358 ( .ip1(n10702), .ip2(\cache_data_A[7][29] ), .op(n12364) );
  nand2_1 U15359 ( .ip1(n12410), .ip2(\cache_data_A[3][29] ), .op(n12363) );
  nand2_1 U15360 ( .ip1(n12242), .ip2(\cache_data_A[1][29] ), .op(n12362) );
  nand2_1 U15361 ( .ip1(n8452), .ip2(\cache_data_A[0][29] ), .op(n12361) );
  nand4_1 U15362 ( .ip1(n12364), .ip2(n12363), .ip3(n12362), .ip4(n12361), 
        .op(n12365) );
  not_ab_or_c_or_d U15363 ( .ip1(\cache_data_A[2][29] ), .ip2(n12546), .ip3(
        n12366), .ip4(n12365), .op(n12368) );
  nand2_1 U15364 ( .ip1(n12582), .ip2(\cache_data_A[5][29] ), .op(n12367) );
  nand3_1 U15365 ( .ip1(n12369), .ip2(n12368), .ip3(n12367), .op(n13128) );
  nand2_1 U15366 ( .ip1(n12550), .ip2(n13128), .op(n12392) );
  nand2_1 U15367 ( .ip1(\cache_data_B[0][93] ), .ip2(n12370), .op(n12380) );
  and2_1 U15368 ( .ip1(n12581), .ip2(\cache_data_B[7][93] ), .op(n12377) );
  nand2_1 U15369 ( .ip1(n11280), .ip2(\cache_data_B[5][93] ), .op(n12375) );
  nand2_1 U15370 ( .ip1(n12371), .ip2(\cache_data_B[6][93] ), .op(n12374) );
  nand2_1 U15371 ( .ip1(n8060), .ip2(\cache_data_B[3][93] ), .op(n12373) );
  nand2_1 U15372 ( .ip1(n11946), .ip2(\cache_data_B[1][93] ), .op(n12372) );
  nand4_1 U15373 ( .ip1(n12375), .ip2(n12374), .ip3(n12373), .ip4(n12372), 
        .op(n12376) );
  not_ab_or_c_or_d U15374 ( .ip1(\cache_data_B[2][93] ), .ip2(n12546), .ip3(
        n12377), .ip4(n12376), .op(n12379) );
  nand2_1 U15375 ( .ip1(n12476), .ip2(\cache_data_B[4][93] ), .op(n12378) );
  nand3_1 U15376 ( .ip1(n12380), .ip2(n12379), .ip3(n12378), .op(n13129) );
  nand2_1 U15377 ( .ip1(n12580), .ip2(n13129), .op(n12391) );
  nand2_1 U15378 ( .ip1(n12429), .ip2(\cache_data_B[6][61] ), .op(n12389) );
  and2_1 U15379 ( .ip1(n12591), .ip2(\cache_data_B[3][61] ), .op(n12386) );
  nand2_1 U15380 ( .ip1(n11304), .ip2(\cache_data_B[5][61] ), .op(n12384) );
  nand2_1 U15381 ( .ip1(n12475), .ip2(\cache_data_B[2][61] ), .op(n12383) );
  nand2_1 U15382 ( .ip1(n12552), .ip2(\cache_data_B[7][61] ), .op(n12382) );
  nand2_1 U15383 ( .ip1(n12396), .ip2(\cache_data_B[4][61] ), .op(n12381) );
  nand4_1 U15384 ( .ip1(n12384), .ip2(n12383), .ip3(n12382), .ip4(n12381), 
        .op(n12385) );
  not_ab_or_c_or_d U15385 ( .ip1(\cache_data_B[0][61] ), .ip2(n12204), .ip3(
        n12386), .ip4(n12385), .op(n12388) );
  nand2_1 U15386 ( .ip1(n11946), .ip2(\cache_data_B[1][61] ), .op(n12387) );
  nand3_1 U15387 ( .ip1(n12389), .ip2(n12388), .ip3(n12387), .op(n13137) );
  nand2_1 U15388 ( .ip1(n12563), .ip2(n13137), .op(n12390) );
  nand4_1 U15389 ( .ip1(n12393), .ip2(n12392), .ip3(n12391), .ip4(n12390), 
        .op(n12394) );
  not_ab_or_c_or_d U15390 ( .ip1(n12509), .ip2(n13130), .ip3(n12395), .ip4(
        n12394), .op(n12407) );
  nand2_1 U15391 ( .ip1(\cache_data_A[6][61] ), .ip2(n12458), .op(n12405) );
  and2_1 U15392 ( .ip1(n12396), .ip2(\cache_data_A[4][61] ), .op(n12402) );
  nand2_1 U15393 ( .ip1(n8060), .ip2(\cache_data_A[3][61] ), .op(n12400) );
  nand2_1 U15394 ( .ip1(n8452), .ip2(\cache_data_A[0][61] ), .op(n12399) );
  nand2_1 U15395 ( .ip1(n10166), .ip2(\cache_data_A[1][61] ), .op(n12398) );
  nand2_1 U15396 ( .ip1(n12581), .ip2(\cache_data_A[7][61] ), .op(n12397) );
  nand4_1 U15397 ( .ip1(n12400), .ip2(n12399), .ip3(n12398), .ip4(n12397), 
        .op(n12401) );
  not_ab_or_c_or_d U15398 ( .ip1(n12546), .ip2(\cache_data_A[2][61] ), .ip3(
        n12402), .ip4(n12401), .op(n12404) );
  nand2_1 U15399 ( .ip1(n12582), .ip2(\cache_data_A[5][61] ), .op(n12403) );
  nand3_1 U15400 ( .ip1(n12405), .ip2(n12404), .ip3(n12403), .op(n13138) );
  nand2_1 U15401 ( .ip1(n12595), .ip2(n13138), .op(n12406) );
  nand3_1 U15402 ( .ip1(n12408), .ip2(n12407), .ip3(n12406), .op(n12409) );
  mux2_1 U15403 ( .ip1(N4117), .ip2(n12409), .s(n12599), .op(n5291) );
  nand2_1 U15404 ( .ip1(\cache_data_A[3][62] ), .ip2(n12410), .op(n12419) );
  and2_1 U15405 ( .ip1(n12256), .ip2(\cache_data_A[5][62] ), .op(n12416) );
  nand2_1 U15406 ( .ip1(n12581), .ip2(\cache_data_A[7][62] ), .op(n12414) );
  nand2_1 U15407 ( .ip1(n12297), .ip2(\cache_data_A[0][62] ), .op(n12413) );
  nand2_1 U15408 ( .ip1(n12475), .ip2(\cache_data_A[2][62] ), .op(n12412) );
  nand2_1 U15409 ( .ip1(n12242), .ip2(\cache_data_A[1][62] ), .op(n12411) );
  nand4_1 U15410 ( .ip1(n12414), .ip2(n12413), .ip3(n12412), .ip4(n12411), 
        .op(n12415) );
  not_ab_or_c_or_d U15411 ( .ip1(n12551), .ip2(\cache_data_A[6][62] ), .ip3(
        n12416), .ip4(n12415), .op(n12418) );
  nand2_1 U15412 ( .ip1(n12476), .ip2(\cache_data_A[4][62] ), .op(n12417) );
  nand3_1 U15413 ( .ip1(n12419), .ip2(n12418), .ip3(n12417), .op(n13143) );
  nand2_1 U15414 ( .ip1(n12595), .ip2(n13143), .op(n12498) );
  nand2_1 U15415 ( .ip1(\cache_data_A[7][126] ), .ip2(n12468), .op(n12428) );
  and2_1 U15416 ( .ip1(n11724), .ip2(\cache_data_A[1][126] ), .op(n12425) );
  nand2_1 U15417 ( .ip1(n12582), .ip2(\cache_data_A[5][126] ), .op(n12423) );
  nand2_1 U15418 ( .ip1(n11855), .ip2(\cache_data_A[2][126] ), .op(n12422) );
  nand2_1 U15419 ( .ip1(n12476), .ip2(\cache_data_A[4][126] ), .op(n12421) );
  nand2_1 U15420 ( .ip1(n12321), .ip2(\cache_data_A[3][126] ), .op(n12420) );
  nand4_1 U15421 ( .ip1(n12423), .ip2(n12422), .ip3(n12421), .ip4(n12420), 
        .op(n12424) );
  not_ab_or_c_or_d U15422 ( .ip1(\cache_data_A[0][126] ), .ip2(n12204), .ip3(
        n12425), .ip4(n12424), .op(n12427) );
  nand2_1 U15423 ( .ip1(n12429), .ip2(\cache_data_A[6][126] ), .op(n12426) );
  nand3_1 U15424 ( .ip1(n12428), .ip2(n12427), .ip3(n12426), .op(n13155) );
  nand2_1 U15425 ( .ip1(n12486), .ip2(\cache_data_A[2][94] ), .op(n12433) );
  nand2_1 U15426 ( .ip1(n11946), .ip2(\cache_data_A[1][94] ), .op(n12432) );
  nand2_1 U15427 ( .ip1(n12429), .ip2(\cache_data_A[6][94] ), .op(n12431) );
  nand2_1 U15428 ( .ip1(n12256), .ip2(\cache_data_A[5][94] ), .op(n12430) );
  nand4_1 U15429 ( .ip1(n12433), .ip2(n12432), .ip3(n12431), .ip4(n12430), 
        .op(n12439) );
  nand2_1 U15430 ( .ip1(n8452), .ip2(\cache_data_A[0][94] ), .op(n12437) );
  nand2_1 U15431 ( .ip1(n12581), .ip2(\cache_data_A[7][94] ), .op(n12436) );
  nand2_1 U15432 ( .ip1(n12321), .ip2(\cache_data_A[3][94] ), .op(n12435) );
  nand2_1 U15433 ( .ip1(n12476), .ip2(\cache_data_A[4][94] ), .op(n12434) );
  nand4_1 U15434 ( .ip1(n12437), .ip2(n12436), .ip3(n12435), .ip4(n12434), 
        .op(n12438) );
  nor2_1 U15435 ( .ip1(n12439), .ip2(n12438), .op(n13144) );
  nor2_1 U15436 ( .ip1(n13144), .ip2(n12529), .op(n12485) );
  nand2_1 U15437 ( .ip1(n12475), .ip2(\cache_data_A[2][30] ), .op(n12448) );
  and2_1 U15438 ( .ip1(n11296), .ip2(\cache_data_A[5][30] ), .op(n12445) );
  nand2_1 U15439 ( .ip1(n8060), .ip2(\cache_data_A[3][30] ), .op(n12443) );
  nand2_1 U15440 ( .ip1(n12581), .ip2(\cache_data_A[7][30] ), .op(n12442) );
  nand2_1 U15441 ( .ip1(n12297), .ip2(\cache_data_A[0][30] ), .op(n12441) );
  nand2_1 U15442 ( .ip1(n10686), .ip2(\cache_data_A[1][30] ), .op(n12440) );
  nand4_1 U15443 ( .ip1(n12443), .ip2(n12442), .ip3(n12441), .ip4(n12440), 
        .op(n12444) );
  not_ab_or_c_or_d U15444 ( .ip1(\cache_data_A[6][30] ), .ip2(n12551), .ip3(
        n12445), .ip4(n12444), .op(n12447) );
  nand2_1 U15445 ( .ip1(n12476), .ip2(\cache_data_A[4][30] ), .op(n12446) );
  nand3_1 U15446 ( .ip1(n12448), .ip2(n12447), .ip3(n12446), .op(n13146) );
  nand2_1 U15447 ( .ip1(n12550), .ip2(n13146), .op(n12483) );
  nand2_1 U15448 ( .ip1(n12476), .ip2(\cache_data_B[4][30] ), .op(n12457) );
  and2_1 U15449 ( .ip1(n12320), .ip2(\cache_data_B[6][30] ), .op(n12454) );
  nand2_1 U15450 ( .ip1(n8060), .ip2(\cache_data_B[3][30] ), .op(n12452) );
  nand2_1 U15451 ( .ip1(n8452), .ip2(\cache_data_B[0][30] ), .op(n12451) );
  nand2_1 U15452 ( .ip1(n12581), .ip2(\cache_data_B[7][30] ), .op(n12450) );
  nand2_1 U15453 ( .ip1(n12582), .ip2(\cache_data_B[5][30] ), .op(n12449) );
  nand4_1 U15454 ( .ip1(n12452), .ip2(n12451), .ip3(n12450), .ip4(n12449), 
        .op(n12453) );
  not_ab_or_c_or_d U15455 ( .ip1(n12546), .ip2(\cache_data_B[2][30] ), .ip3(
        n12454), .ip4(n12453), .op(n12456) );
  nand2_1 U15456 ( .ip1(n12242), .ip2(\cache_data_B[1][30] ), .op(n12455) );
  nand3_1 U15457 ( .ip1(n12457), .ip2(n12456), .ip3(n12455), .op(n13148) );
  nand2_1 U15458 ( .ip1(n12539), .ip2(n13148), .op(n12482) );
  nand2_1 U15459 ( .ip1(\cache_data_B[3][126] ), .ip2(n8060), .op(n12467) );
  and2_1 U15460 ( .ip1(n12582), .ip2(\cache_data_B[5][126] ), .op(n12464) );
  nand2_1 U15461 ( .ip1(n10702), .ip2(\cache_data_B[7][126] ), .op(n12462) );
  nand2_1 U15462 ( .ip1(n12458), .ip2(\cache_data_B[6][126] ), .op(n12461) );
  nand2_1 U15463 ( .ip1(n12475), .ip2(\cache_data_B[2][126] ), .op(n12460) );
  nand2_1 U15464 ( .ip1(n8452), .ip2(\cache_data_B[0][126] ), .op(n12459) );
  nand4_1 U15465 ( .ip1(n12462), .ip2(n12461), .ip3(n12460), .ip4(n12459), 
        .op(n12463) );
  not_ab_or_c_or_d U15466 ( .ip1(n11324), .ip2(\cache_data_B[4][126] ), .ip3(
        n12464), .ip4(n12463), .op(n12466) );
  nand2_1 U15467 ( .ip1(n11311), .ip2(\cache_data_B[1][126] ), .op(n12465) );
  nand3_1 U15468 ( .ip1(n12467), .ip2(n12466), .ip3(n12465), .op(n13145) );
  nand2_1 U15469 ( .ip1(n12573), .ip2(n13145), .op(n12481) );
  nand2_1 U15470 ( .ip1(n12468), .ip2(\cache_data_B[7][94] ), .op(n12479) );
  and2_1 U15471 ( .ip1(n10686), .ip2(\cache_data_B[1][94] ), .op(n12474) );
  nand2_1 U15472 ( .ip1(n12321), .ip2(\cache_data_B[3][94] ), .op(n12472) );
  nand2_1 U15473 ( .ip1(n12582), .ip2(\cache_data_B[5][94] ), .op(n12471) );
  nand2_1 U15474 ( .ip1(n12297), .ip2(\cache_data_B[0][94] ), .op(n12470) );
  nand2_1 U15475 ( .ip1(n12551), .ip2(\cache_data_B[6][94] ), .op(n12469) );
  nand4_1 U15476 ( .ip1(n12472), .ip2(n12471), .ip3(n12470), .ip4(n12469), 
        .op(n12473) );
  not_ab_or_c_or_d U15477 ( .ip1(\cache_data_B[2][94] ), .ip2(n12475), .ip3(
        n12474), .ip4(n12473), .op(n12478) );
  nand2_1 U15478 ( .ip1(n12476), .ip2(\cache_data_B[4][94] ), .op(n12477) );
  nand3_1 U15479 ( .ip1(n12479), .ip2(n12478), .ip3(n12477), .op(n13147) );
  nand2_1 U15480 ( .ip1(n12580), .ip2(n13147), .op(n12480) );
  nand4_1 U15481 ( .ip1(n12483), .ip2(n12482), .ip3(n12481), .ip4(n12480), 
        .op(n12484) );
  not_ab_or_c_or_d U15482 ( .ip1(n12509), .ip2(n13155), .ip3(n12485), .ip4(
        n12484), .op(n12497) );
  nand2_1 U15483 ( .ip1(\cache_data_B[2][62] ), .ip2(n12486), .op(n12495) );
  and2_1 U15484 ( .ip1(n10166), .ip2(\cache_data_B[1][62] ), .op(n12492) );
  nand2_1 U15485 ( .ip1(n12584), .ip2(\cache_data_B[4][62] ), .op(n12490) );
  nand2_1 U15486 ( .ip1(n12551), .ip2(\cache_data_B[6][62] ), .op(n12489) );
  nand2_1 U15487 ( .ip1(n8452), .ip2(\cache_data_B[0][62] ), .op(n12488) );
  nand2_1 U15488 ( .ip1(n12581), .ip2(\cache_data_B[7][62] ), .op(n12487) );
  nand4_1 U15489 ( .ip1(n12490), .ip2(n12489), .ip3(n12488), .ip4(n12487), 
        .op(n12491) );
  not_ab_or_c_or_d U15490 ( .ip1(\cache_data_B[3][62] ), .ip2(n12559), .ip3(
        n12492), .ip4(n12491), .op(n12494) );
  nand2_1 U15491 ( .ip1(n12118), .ip2(\cache_data_B[5][62] ), .op(n12493) );
  nand3_1 U15492 ( .ip1(n12495), .ip2(n12494), .ip3(n12493), .op(n13156) );
  nand2_1 U15493 ( .ip1(n12563), .ip2(n13156), .op(n12496) );
  nand3_1 U15494 ( .ip1(n12498), .ip2(n12497), .ip3(n12496), .op(n12499) );
  mux2_1 U15495 ( .ip1(N4114), .ip2(n12499), .s(n12599), .op(n5290) );
  nand2_1 U15496 ( .ip1(n11142), .ip2(\cache_data_A[2][127] ), .op(n12508) );
  and2_1 U15497 ( .ip1(n12584), .ip2(\cache_data_A[4][127] ), .op(n12505) );
  nand2_1 U15498 ( .ip1(n11311), .ip2(\cache_data_A[1][127] ), .op(n12503) );
  nand2_1 U15499 ( .ip1(n12551), .ip2(\cache_data_A[6][127] ), .op(n12502) );
  nand2_1 U15500 ( .ip1(n11057), .ip2(\cache_data_A[7][127] ), .op(n12501) );
  nand2_1 U15501 ( .ip1(n12204), .ip2(\cache_data_A[0][127] ), .op(n12500) );
  nand4_1 U15502 ( .ip1(n12503), .ip2(n12502), .ip3(n12501), .ip4(n12500), 
        .op(n12504) );
  not_ab_or_c_or_d U15503 ( .ip1(\cache_data_A[3][127] ), .ip2(n12559), .ip3(
        n12505), .ip4(n12504), .op(n12507) );
  nand2_1 U15504 ( .ip1(n12582), .ip2(\cache_data_A[5][127] ), .op(n12506) );
  nand3_1 U15505 ( .ip1(n12508), .ip2(n12507), .ip3(n12506), .op(n13171) );
  nand2_1 U15506 ( .ip1(n12509), .ip2(n13171), .op(n12598) );
  nand2_1 U15507 ( .ip1(n12584), .ip2(\cache_data_B[4][95] ), .op(n12518) );
  and2_1 U15508 ( .ip1(n12581), .ip2(\cache_data_B[7][95] ), .op(n12515) );
  nand2_1 U15509 ( .ip1(n12559), .ip2(\cache_data_B[3][95] ), .op(n12513) );
  nand2_1 U15510 ( .ip1(n12551), .ip2(\cache_data_B[6][95] ), .op(n12512) );
  nand2_1 U15511 ( .ip1(n11946), .ip2(\cache_data_B[1][95] ), .op(n12511) );
  nand2_1 U15512 ( .ip1(n12583), .ip2(\cache_data_B[2][95] ), .op(n12510) );
  nand4_1 U15513 ( .ip1(n12513), .ip2(n12512), .ip3(n12511), .ip4(n12510), 
        .op(n12514) );
  not_ab_or_c_or_d U15514 ( .ip1(n11911), .ip2(\cache_data_B[0][95] ), .ip3(
        n12515), .ip4(n12514), .op(n12517) );
  nand2_1 U15515 ( .ip1(n12582), .ip2(\cache_data_B[5][95] ), .op(n12516) );
  nand3_1 U15516 ( .ip1(n12518), .ip2(n12517), .ip3(n12516), .op(n13167) );
  nand2_1 U15517 ( .ip1(n12583), .ip2(\cache_data_A[2][95] ), .op(n12522) );
  nand2_1 U15518 ( .ip1(n12581), .ip2(\cache_data_A[7][95] ), .op(n12521) );
  nand2_1 U15519 ( .ip1(n8060), .ip2(\cache_data_A[3][95] ), .op(n12520) );
  nand2_1 U15520 ( .ip1(n12582), .ip2(\cache_data_A[5][95] ), .op(n12519) );
  nand4_1 U15521 ( .ip1(n12522), .ip2(n12521), .ip3(n12520), .ip4(n12519), 
        .op(n12528) );
  nand2_1 U15522 ( .ip1(n12584), .ip2(\cache_data_A[4][95] ), .op(n12526) );
  nand2_1 U15523 ( .ip1(n10686), .ip2(\cache_data_A[1][95] ), .op(n12525) );
  nand2_1 U15524 ( .ip1(n12551), .ip2(\cache_data_A[6][95] ), .op(n12524) );
  nand2_1 U15525 ( .ip1(n12297), .ip2(\cache_data_A[0][95] ), .op(n12523) );
  nand4_1 U15526 ( .ip1(n12526), .ip2(n12525), .ip3(n12524), .ip4(n12523), 
        .op(n12527) );
  nor2_1 U15527 ( .ip1(n12528), .ip2(n12527), .op(n13164) );
  nor2_1 U15528 ( .ip1(n13164), .ip2(n12529), .op(n12579) );
  nand2_1 U15529 ( .ip1(n12551), .ip2(\cache_data_B[6][31] ), .op(n12538) );
  and2_1 U15530 ( .ip1(n11304), .ip2(\cache_data_B[5][31] ), .op(n12535) );
  nand2_1 U15531 ( .ip1(n12581), .ip2(\cache_data_B[7][31] ), .op(n12533) );
  nand2_1 U15532 ( .ip1(n12584), .ip2(\cache_data_B[4][31] ), .op(n12532) );
  nand2_1 U15533 ( .ip1(n12297), .ip2(\cache_data_B[0][31] ), .op(n12531) );
  nand2_1 U15534 ( .ip1(n11946), .ip2(\cache_data_B[1][31] ), .op(n12530) );
  nand4_1 U15535 ( .ip1(n12533), .ip2(n12532), .ip3(n12531), .ip4(n12530), 
        .op(n12534) );
  not_ab_or_c_or_d U15536 ( .ip1(n12546), .ip2(\cache_data_B[2][31] ), .ip3(
        n12535), .ip4(n12534), .op(n12537) );
  nand2_1 U15537 ( .ip1(n12321), .ip2(\cache_data_B[3][31] ), .op(n12536) );
  nand3_1 U15538 ( .ip1(n12538), .ip2(n12537), .ip3(n12536), .op(n13169) );
  nand2_1 U15539 ( .ip1(n12539), .ip2(n13169), .op(n12577) );
  nand2_1 U15540 ( .ip1(n12357), .ip2(\cache_data_A[0][31] ), .op(n12549) );
  and2_1 U15541 ( .ip1(n11780), .ip2(\cache_data_A[6][31] ), .op(n12545) );
  nand2_1 U15542 ( .ip1(n12581), .ip2(\cache_data_A[7][31] ), .op(n12543) );
  nand2_1 U15543 ( .ip1(n12321), .ip2(\cache_data_A[3][31] ), .op(n12542) );
  nand2_1 U15544 ( .ip1(n11311), .ip2(\cache_data_A[1][31] ), .op(n12541) );
  nand2_1 U15545 ( .ip1(n12582), .ip2(\cache_data_A[5][31] ), .op(n12540) );
  nand4_1 U15546 ( .ip1(n12543), .ip2(n12542), .ip3(n12541), .ip4(n12540), 
        .op(n12544) );
  not_ab_or_c_or_d U15547 ( .ip1(\cache_data_A[2][31] ), .ip2(n12546), .ip3(
        n12545), .ip4(n12544), .op(n12548) );
  nand2_1 U15548 ( .ip1(n12584), .ip2(\cache_data_A[4][31] ), .op(n12547) );
  nand3_1 U15549 ( .ip1(n12549), .ip2(n12548), .ip3(n12547), .op(n13179) );
  nand2_1 U15550 ( .ip1(n12550), .ip2(n13179), .op(n12576) );
  nand2_1 U15551 ( .ip1(n12551), .ip2(\cache_data_B[6][63] ), .op(n12562) );
  and2_1 U15552 ( .ip1(n12476), .ip2(\cache_data_B[4][63] ), .op(n12558) );
  nand2_1 U15553 ( .ip1(n12552), .ip2(\cache_data_B[7][63] ), .op(n12556) );
  nand2_1 U15554 ( .ip1(n12583), .ip2(\cache_data_B[2][63] ), .op(n12555) );
  nand2_1 U15555 ( .ip1(n12582), .ip2(\cache_data_B[5][63] ), .op(n12554) );
  nand2_1 U15556 ( .ip1(n12297), .ip2(\cache_data_B[0][63] ), .op(n12553) );
  nand4_1 U15557 ( .ip1(n12556), .ip2(n12555), .ip3(n12554), .ip4(n12553), 
        .op(n12557) );
  not_ab_or_c_or_d U15558 ( .ip1(\cache_data_B[3][63] ), .ip2(n12559), .ip3(
        n12558), .ip4(n12557), .op(n12561) );
  nand2_1 U15559 ( .ip1(n11946), .ip2(\cache_data_B[1][63] ), .op(n12560) );
  nand3_1 U15560 ( .ip1(n12562), .ip2(n12561), .ip3(n12560), .op(n13181) );
  nand2_1 U15561 ( .ip1(n12563), .ip2(n13181), .op(n12575) );
  nand2_1 U15562 ( .ip1(n12584), .ip2(\cache_data_B[4][127] ), .op(n12572) );
  and2_1 U15563 ( .ip1(n12429), .ip2(\cache_data_B[6][127] ), .op(n12569) );
  nand2_1 U15564 ( .ip1(n8060), .ip2(\cache_data_B[3][127] ), .op(n12567) );
  nand2_1 U15565 ( .ip1(n10686), .ip2(\cache_data_B[1][127] ), .op(n12566) );
  nand2_1 U15566 ( .ip1(n12581), .ip2(\cache_data_B[7][127] ), .op(n12565) );
  nand2_1 U15567 ( .ip1(n12583), .ip2(\cache_data_B[2][127] ), .op(n12564) );
  nand4_1 U15568 ( .ip1(n12567), .ip2(n12566), .ip3(n12565), .ip4(n12564), 
        .op(n12568) );
  not_ab_or_c_or_d U15569 ( .ip1(n11911), .ip2(\cache_data_B[0][127] ), .ip3(
        n12569), .ip4(n12568), .op(n12571) );
  nand2_1 U15570 ( .ip1(n12582), .ip2(\cache_data_B[5][127] ), .op(n12570) );
  nand3_1 U15571 ( .ip1(n12572), .ip2(n12571), .ip3(n12570), .op(n13165) );
  nand2_1 U15572 ( .ip1(n12573), .ip2(n13165), .op(n12574) );
  nand4_1 U15573 ( .ip1(n12577), .ip2(n12576), .ip3(n12575), .ip4(n12574), 
        .op(n12578) );
  not_ab_or_c_or_d U15574 ( .ip1(n12580), .ip2(n13167), .ip3(n12579), .ip4(
        n12578), .op(n12597) );
  nand2_1 U15575 ( .ip1(n12581), .ip2(\cache_data_A[7][63] ), .op(n12594) );
  and2_1 U15576 ( .ip1(n12371), .ip2(\cache_data_A[6][63] ), .op(n12590) );
  nand2_1 U15577 ( .ip1(n12582), .ip2(\cache_data_A[5][63] ), .op(n12588) );
  nand2_1 U15578 ( .ip1(n11311), .ip2(\cache_data_A[1][63] ), .op(n12587) );
  nand2_1 U15579 ( .ip1(n12583), .ip2(\cache_data_A[2][63] ), .op(n12586) );
  nand2_1 U15580 ( .ip1(n12584), .ip2(\cache_data_A[4][63] ), .op(n12585) );
  nand4_1 U15581 ( .ip1(n12588), .ip2(n12587), .ip3(n12586), .ip4(n12585), 
        .op(n12589) );
  not_ab_or_c_or_d U15582 ( .ip1(n8452), .ip2(\cache_data_A[0][63] ), .ip3(
        n12590), .ip4(n12589), .op(n12593) );
  nand2_1 U15583 ( .ip1(n12591), .ip2(\cache_data_A[3][63] ), .op(n12592) );
  nand3_1 U15584 ( .ip1(n12594), .ip2(n12593), .ip3(n12592), .op(n13161) );
  nand2_1 U15585 ( .ip1(n12595), .ip2(n13161), .op(n12596) );
  nand3_1 U15586 ( .ip1(n12598), .ip2(n12597), .ip3(n12596), .op(n12600) );
  mux2_1 U15587 ( .ip1(N4111), .ip2(n12600), .s(n12599), .op(n5289) );
  nand2_1 U15588 ( .ip1(n13172), .ip2(n12601), .op(n12617) );
  nor2_1 U15589 ( .ip1(n12602), .ip2(n13163), .op(n12612) );
  nand2_1 U15590 ( .ip1(n13168), .ip2(n12603), .op(n12610) );
  nand2_1 U15591 ( .ip1(n13162), .ip2(n12604), .op(n12609) );
  nand2_1 U15592 ( .ip1(n13180), .ip2(n12605), .op(n12608) );
  nand2_1 U15593 ( .ip1(n13166), .ip2(n12606), .op(n12607) );
  nand4_1 U15594 ( .ip1(n12610), .ip2(n12609), .ip3(n12608), .ip4(n12607), 
        .op(n12611) );
  not_ab_or_c_or_d U15595 ( .ip1(n13170), .ip2(n12613), .ip3(n12612), .ip4(
        n12611), .op(n12616) );
  nand2_1 U15596 ( .ip1(n13182), .ip2(n12614), .op(n12615) );
  nand3_1 U15597 ( .ip1(n12617), .ip2(n12616), .ip3(n12615), .op(n12619) );
  nor2_1 U15598 ( .ip1(n12618), .ip2(n13189), .op(n13033) );
  mux2_1 U15599 ( .ip1(data_wr_mem[0]), .ip2(n12619), .s(n13033), .op(n5288)
         );
  nand2_1 U15600 ( .ip1(n13172), .ip2(n12620), .op(n12636) );
  nor2_1 U15601 ( .ip1(n12621), .ip2(n13163), .op(n12631) );
  nand2_1 U15602 ( .ip1(n13162), .ip2(n12622), .op(n12629) );
  nand2_1 U15603 ( .ip1(n13180), .ip2(n12623), .op(n12628) );
  nand2_1 U15604 ( .ip1(n13166), .ip2(n12624), .op(n12627) );
  nand2_1 U15605 ( .ip1(n13182), .ip2(n12625), .op(n12626) );
  nand4_1 U15606 ( .ip1(n12629), .ip2(n12628), .ip3(n12627), .ip4(n12626), 
        .op(n12630) );
  not_ab_or_c_or_d U15607 ( .ip1(n13168), .ip2(n12632), .ip3(n12631), .ip4(
        n12630), .op(n12635) );
  nand2_1 U15608 ( .ip1(n13170), .ip2(n12633), .op(n12634) );
  nand3_1 U15609 ( .ip1(n12636), .ip2(n12635), .ip3(n12634), .op(n12637) );
  mux2_1 U15610 ( .ip1(data_wr_mem[1]), .ip2(n12637), .s(n13033), .op(n5287)
         );
  nand2_1 U15611 ( .ip1(n13180), .ip2(n12638), .op(n12654) );
  nor2_1 U15612 ( .ip1(n12639), .ip2(n13163), .op(n12649) );
  nand2_1 U15613 ( .ip1(n13168), .ip2(n12640), .op(n12647) );
  nand2_1 U15614 ( .ip1(n13170), .ip2(n12641), .op(n12646) );
  nand2_1 U15615 ( .ip1(n13166), .ip2(n12642), .op(n12645) );
  nand2_1 U15616 ( .ip1(n13182), .ip2(n12643), .op(n12644) );
  nand4_1 U15617 ( .ip1(n12647), .ip2(n12646), .ip3(n12645), .ip4(n12644), 
        .op(n12648) );
  not_ab_or_c_or_d U15618 ( .ip1(n13172), .ip2(n12650), .ip3(n12649), .ip4(
        n12648), .op(n12653) );
  nand2_1 U15619 ( .ip1(n13162), .ip2(n12651), .op(n12652) );
  nand3_1 U15620 ( .ip1(n12654), .ip2(n12653), .ip3(n12652), .op(n12655) );
  mux2_1 U15621 ( .ip1(data_wr_mem[2]), .ip2(n12655), .s(n13033), .op(n5286)
         );
  nand2_1 U15622 ( .ip1(n13172), .ip2(n12656), .op(n12672) );
  nor2_1 U15623 ( .ip1(n12657), .ip2(n13163), .op(n12667) );
  nand2_1 U15624 ( .ip1(n13166), .ip2(n12658), .op(n12665) );
  nand2_1 U15625 ( .ip1(n13170), .ip2(n12659), .op(n12664) );
  nand2_1 U15626 ( .ip1(n13162), .ip2(n12660), .op(n12663) );
  nand2_1 U15627 ( .ip1(n13168), .ip2(n12661), .op(n12662) );
  nand4_1 U15628 ( .ip1(n12665), .ip2(n12664), .ip3(n12663), .ip4(n12662), 
        .op(n12666) );
  not_ab_or_c_or_d U15629 ( .ip1(n13180), .ip2(n12668), .ip3(n12667), .ip4(
        n12666), .op(n12671) );
  nand2_1 U15630 ( .ip1(n13182), .ip2(n12669), .op(n12670) );
  nand3_1 U15631 ( .ip1(n12672), .ip2(n12671), .ip3(n12670), .op(n12673) );
  mux2_1 U15632 ( .ip1(data_wr_mem[3]), .ip2(n12673), .s(n13033), .op(n5285)
         );
  nand2_1 U15633 ( .ip1(n13180), .ip2(n12674), .op(n12690) );
  nor2_1 U15634 ( .ip1(n12675), .ip2(n13163), .op(n12685) );
  nand2_1 U15635 ( .ip1(n13166), .ip2(n12676), .op(n12683) );
  nand2_1 U15636 ( .ip1(n13172), .ip2(n12677), .op(n12682) );
  nand2_1 U15637 ( .ip1(n13182), .ip2(n12678), .op(n12681) );
  nand2_1 U15638 ( .ip1(n13170), .ip2(n12679), .op(n12680) );
  nand4_1 U15639 ( .ip1(n12683), .ip2(n12682), .ip3(n12681), .ip4(n12680), 
        .op(n12684) );
  not_ab_or_c_or_d U15640 ( .ip1(n13168), .ip2(n12686), .ip3(n12685), .ip4(
        n12684), .op(n12689) );
  nand2_1 U15641 ( .ip1(n13162), .ip2(n12687), .op(n12688) );
  nand3_1 U15642 ( .ip1(n12690), .ip2(n12689), .ip3(n12688), .op(n12691) );
  mux2_1 U15643 ( .ip1(data_wr_mem[4]), .ip2(n12691), .s(n13033), .op(n5284)
         );
  nand2_1 U15644 ( .ip1(n13180), .ip2(n12692), .op(n12708) );
  nor2_1 U15645 ( .ip1(n12693), .ip2(n13163), .op(n12703) );
  nand2_1 U15646 ( .ip1(n13166), .ip2(n12694), .op(n12701) );
  nand2_1 U15647 ( .ip1(n13170), .ip2(n12695), .op(n12700) );
  nand2_1 U15648 ( .ip1(n13168), .ip2(n12696), .op(n12699) );
  nand2_1 U15649 ( .ip1(n13182), .ip2(n12697), .op(n12698) );
  nand4_1 U15650 ( .ip1(n12701), .ip2(n12700), .ip3(n12699), .ip4(n12698), 
        .op(n12702) );
  not_ab_or_c_or_d U15651 ( .ip1(n13172), .ip2(n12704), .ip3(n12703), .ip4(
        n12702), .op(n12707) );
  nand2_1 U15652 ( .ip1(n13162), .ip2(n12705), .op(n12706) );
  nand3_1 U15653 ( .ip1(n12708), .ip2(n12707), .ip3(n12706), .op(n12709) );
  mux2_1 U15654 ( .ip1(data_wr_mem[5]), .ip2(n12709), .s(n13033), .op(n5283)
         );
  nand2_1 U15655 ( .ip1(n13180), .ip2(n12710), .op(n12726) );
  nor2_1 U15656 ( .ip1(n12711), .ip2(n13163), .op(n12721) );
  nand2_1 U15657 ( .ip1(n13166), .ip2(n12712), .op(n12719) );
  nand2_1 U15658 ( .ip1(n13168), .ip2(n12713), .op(n12718) );
  nand2_1 U15659 ( .ip1(n13172), .ip2(n12714), .op(n12717) );
  nand2_1 U15660 ( .ip1(n13182), .ip2(n12715), .op(n12716) );
  nand4_1 U15661 ( .ip1(n12719), .ip2(n12718), .ip3(n12717), .ip4(n12716), 
        .op(n12720) );
  not_ab_or_c_or_d U15662 ( .ip1(n13170), .ip2(n12722), .ip3(n12721), .ip4(
        n12720), .op(n12725) );
  nand2_1 U15663 ( .ip1(n13162), .ip2(n12723), .op(n12724) );
  nand3_1 U15664 ( .ip1(n12726), .ip2(n12725), .ip3(n12724), .op(n12727) );
  mux2_1 U15665 ( .ip1(data_wr_mem[6]), .ip2(n12727), .s(n13033), .op(n5282)
         );
  nand2_1 U15666 ( .ip1(n13180), .ip2(n12728), .op(n12744) );
  nor2_1 U15667 ( .ip1(n12729), .ip2(n13163), .op(n12739) );
  nand2_1 U15668 ( .ip1(n13170), .ip2(n12730), .op(n12737) );
  nand2_1 U15669 ( .ip1(n13182), .ip2(n12731), .op(n12736) );
  nand2_1 U15670 ( .ip1(n13162), .ip2(n12732), .op(n12735) );
  nand2_1 U15671 ( .ip1(n13166), .ip2(n12733), .op(n12734) );
  nand4_1 U15672 ( .ip1(n12737), .ip2(n12736), .ip3(n12735), .ip4(n12734), 
        .op(n12738) );
  not_ab_or_c_or_d U15673 ( .ip1(n13172), .ip2(n12740), .ip3(n12739), .ip4(
        n12738), .op(n12743) );
  nand2_1 U15674 ( .ip1(n13168), .ip2(n12741), .op(n12742) );
  nand3_1 U15675 ( .ip1(n12744), .ip2(n12743), .ip3(n12742), .op(n12745) );
  mux2_1 U15676 ( .ip1(data_wr_mem[7]), .ip2(n12745), .s(n13033), .op(n5281)
         );
  nand2_1 U15677 ( .ip1(n13170), .ip2(n12746), .op(n12762) );
  nor2_1 U15678 ( .ip1(n12747), .ip2(n13163), .op(n12757) );
  nand2_1 U15679 ( .ip1(n13172), .ip2(n12748), .op(n12755) );
  nand2_1 U15680 ( .ip1(n13180), .ip2(n12749), .op(n12754) );
  nand2_1 U15681 ( .ip1(n13162), .ip2(n12750), .op(n12753) );
  nand2_1 U15682 ( .ip1(n13168), .ip2(n12751), .op(n12752) );
  nand4_1 U15683 ( .ip1(n12755), .ip2(n12754), .ip3(n12753), .ip4(n12752), 
        .op(n12756) );
  not_ab_or_c_or_d U15684 ( .ip1(n13166), .ip2(n12758), .ip3(n12757), .ip4(
        n12756), .op(n12761) );
  nand2_1 U15685 ( .ip1(n13182), .ip2(n12759), .op(n12760) );
  nand3_1 U15686 ( .ip1(n12762), .ip2(n12761), .ip3(n12760), .op(n12763) );
  mux2_1 U15687 ( .ip1(data_wr_mem[8]), .ip2(n12763), .s(n13033), .op(n5280)
         );
  nand2_1 U15688 ( .ip1(n13180), .ip2(n12764), .op(n12780) );
  nor2_1 U15689 ( .ip1(n12765), .ip2(n13163), .op(n12775) );
  nand2_1 U15690 ( .ip1(n13182), .ip2(n12766), .op(n12773) );
  nand2_1 U15691 ( .ip1(n13162), .ip2(n12767), .op(n12772) );
  nand2_1 U15692 ( .ip1(n13170), .ip2(n12768), .op(n12771) );
  nand2_1 U15693 ( .ip1(n13168), .ip2(n12769), .op(n12770) );
  nand4_1 U15694 ( .ip1(n12773), .ip2(n12772), .ip3(n12771), .ip4(n12770), 
        .op(n12774) );
  not_ab_or_c_or_d U15695 ( .ip1(n13166), .ip2(n12776), .ip3(n12775), .ip4(
        n12774), .op(n12779) );
  nand2_1 U15696 ( .ip1(n13172), .ip2(n12777), .op(n12778) );
  nand3_1 U15697 ( .ip1(n12780), .ip2(n12779), .ip3(n12778), .op(n12781) );
  buf_1 U15698 ( .ip(n13033), .op(n13186) );
  mux2_1 U15699 ( .ip1(data_wr_mem[9]), .ip2(n12781), .s(n13186), .op(n5279)
         );
  nand2_1 U15700 ( .ip1(n13170), .ip2(n12782), .op(n12798) );
  nor2_1 U15701 ( .ip1(n12783), .ip2(n13163), .op(n12793) );
  nand2_1 U15702 ( .ip1(n13172), .ip2(n12784), .op(n12791) );
  nand2_1 U15703 ( .ip1(n13180), .ip2(n12785), .op(n12790) );
  nand2_1 U15704 ( .ip1(n13166), .ip2(n12786), .op(n12789) );
  nand2_1 U15705 ( .ip1(n13182), .ip2(n12787), .op(n12788) );
  nand4_1 U15706 ( .ip1(n12791), .ip2(n12790), .ip3(n12789), .ip4(n12788), 
        .op(n12792) );
  not_ab_or_c_or_d U15707 ( .ip1(n13168), .ip2(n12794), .ip3(n12793), .ip4(
        n12792), .op(n12797) );
  nand2_1 U15708 ( .ip1(n13162), .ip2(n12795), .op(n12796) );
  nand3_1 U15709 ( .ip1(n12798), .ip2(n12797), .ip3(n12796), .op(n12799) );
  mux2_1 U15710 ( .ip1(data_wr_mem[10]), .ip2(n12799), .s(n13186), .op(n5278)
         );
  nand2_1 U15711 ( .ip1(n13168), .ip2(n12800), .op(n12816) );
  nor2_1 U15712 ( .ip1(n12801), .ip2(n13163), .op(n12811) );
  nand2_1 U15713 ( .ip1(n13162), .ip2(n12802), .op(n12809) );
  nand2_1 U15714 ( .ip1(n13180), .ip2(n12803), .op(n12808) );
  nand2_1 U15715 ( .ip1(n13170), .ip2(n12804), .op(n12807) );
  nand2_1 U15716 ( .ip1(n13172), .ip2(n12805), .op(n12806) );
  nand4_1 U15717 ( .ip1(n12809), .ip2(n12808), .ip3(n12807), .ip4(n12806), 
        .op(n12810) );
  not_ab_or_c_or_d U15718 ( .ip1(n13182), .ip2(n12812), .ip3(n12811), .ip4(
        n12810), .op(n12815) );
  nand2_1 U15719 ( .ip1(n13166), .ip2(n12813), .op(n12814) );
  nand3_1 U15720 ( .ip1(n12816), .ip2(n12815), .ip3(n12814), .op(n12817) );
  mux2_1 U15721 ( .ip1(data_wr_mem[11]), .ip2(n12817), .s(n13033), .op(n5277)
         );
  nand2_1 U15722 ( .ip1(n13166), .ip2(n12818), .op(n12834) );
  nor2_1 U15723 ( .ip1(n12819), .ip2(n13163), .op(n12829) );
  nand2_1 U15724 ( .ip1(n13168), .ip2(n12820), .op(n12827) );
  nand2_1 U15725 ( .ip1(n13182), .ip2(n12821), .op(n12826) );
  nand2_1 U15726 ( .ip1(n13172), .ip2(n12822), .op(n12825) );
  nand2_1 U15727 ( .ip1(n13170), .ip2(n12823), .op(n12824) );
  nand4_1 U15728 ( .ip1(n12827), .ip2(n12826), .ip3(n12825), .ip4(n12824), 
        .op(n12828) );
  not_ab_or_c_or_d U15729 ( .ip1(n13180), .ip2(n12830), .ip3(n12829), .ip4(
        n12828), .op(n12833) );
  nand2_1 U15730 ( .ip1(n13162), .ip2(n12831), .op(n12832) );
  nand3_1 U15731 ( .ip1(n12834), .ip2(n12833), .ip3(n12832), .op(n12835) );
  mux2_1 U15732 ( .ip1(data_wr_mem[12]), .ip2(n12835), .s(n13033), .op(n5276)
         );
  nand2_1 U15733 ( .ip1(n13162), .ip2(n12836), .op(n12852) );
  nor2_1 U15734 ( .ip1(n12837), .ip2(n13163), .op(n12847) );
  nand2_1 U15735 ( .ip1(n13172), .ip2(n12838), .op(n12845) );
  nand2_1 U15736 ( .ip1(n13170), .ip2(n12839), .op(n12844) );
  nand2_1 U15737 ( .ip1(n13168), .ip2(n12840), .op(n12843) );
  nand2_1 U15738 ( .ip1(n13182), .ip2(n12841), .op(n12842) );
  nand4_1 U15739 ( .ip1(n12845), .ip2(n12844), .ip3(n12843), .ip4(n12842), 
        .op(n12846) );
  not_ab_or_c_or_d U15740 ( .ip1(n13180), .ip2(n12848), .ip3(n12847), .ip4(
        n12846), .op(n12851) );
  nand2_1 U15741 ( .ip1(n13166), .ip2(n12849), .op(n12850) );
  nand3_1 U15742 ( .ip1(n12852), .ip2(n12851), .ip3(n12850), .op(n12853) );
  mux2_1 U15743 ( .ip1(data_wr_mem[13]), .ip2(n12853), .s(n13186), .op(n5275)
         );
  nand2_1 U15744 ( .ip1(n13172), .ip2(n12854), .op(n12870) );
  nor2_1 U15745 ( .ip1(n12855), .ip2(n13163), .op(n12865) );
  nand2_1 U15746 ( .ip1(n13180), .ip2(n12856), .op(n12863) );
  nand2_1 U15747 ( .ip1(n13168), .ip2(n12857), .op(n12862) );
  nand2_1 U15748 ( .ip1(n13170), .ip2(n12858), .op(n12861) );
  nand2_1 U15749 ( .ip1(n13182), .ip2(n12859), .op(n12860) );
  nand4_1 U15750 ( .ip1(n12863), .ip2(n12862), .ip3(n12861), .ip4(n12860), 
        .op(n12864) );
  not_ab_or_c_or_d U15751 ( .ip1(n13166), .ip2(n12866), .ip3(n12865), .ip4(
        n12864), .op(n12869) );
  nand2_1 U15752 ( .ip1(n13162), .ip2(n12867), .op(n12868) );
  nand3_1 U15753 ( .ip1(n12870), .ip2(n12869), .ip3(n12868), .op(n12871) );
  mux2_1 U15754 ( .ip1(data_wr_mem[14]), .ip2(n12871), .s(n13033), .op(n5274)
         );
  nand2_1 U15755 ( .ip1(n13172), .ip2(n12872), .op(n12888) );
  nor2_1 U15756 ( .ip1(n12873), .ip2(n13163), .op(n12883) );
  nand2_1 U15757 ( .ip1(n13166), .ip2(n12874), .op(n12881) );
  nand2_1 U15758 ( .ip1(n13182), .ip2(n12875), .op(n12880) );
  nand2_1 U15759 ( .ip1(n13168), .ip2(n12876), .op(n12879) );
  nand2_1 U15760 ( .ip1(n13170), .ip2(n12877), .op(n12878) );
  nand4_1 U15761 ( .ip1(n12881), .ip2(n12880), .ip3(n12879), .ip4(n12878), 
        .op(n12882) );
  not_ab_or_c_or_d U15762 ( .ip1(n13180), .ip2(n12884), .ip3(n12883), .ip4(
        n12882), .op(n12887) );
  nand2_1 U15763 ( .ip1(n13162), .ip2(n12885), .op(n12886) );
  nand3_1 U15764 ( .ip1(n12888), .ip2(n12887), .ip3(n12886), .op(n12889) );
  mux2_1 U15765 ( .ip1(data_wr_mem[15]), .ip2(n12889), .s(n13033), .op(n5273)
         );
  nand2_1 U15766 ( .ip1(n13168), .ip2(n12890), .op(n12906) );
  nor2_1 U15767 ( .ip1(n12891), .ip2(n13163), .op(n12901) );
  nand2_1 U15768 ( .ip1(n13170), .ip2(n12892), .op(n12899) );
  nand2_1 U15769 ( .ip1(n13182), .ip2(n12893), .op(n12898) );
  nand2_1 U15770 ( .ip1(n13162), .ip2(n12894), .op(n12897) );
  nand2_1 U15771 ( .ip1(n13172), .ip2(n12895), .op(n12896) );
  nand4_1 U15772 ( .ip1(n12899), .ip2(n12898), .ip3(n12897), .ip4(n12896), 
        .op(n12900) );
  not_ab_or_c_or_d U15773 ( .ip1(n13180), .ip2(n12902), .ip3(n12901), .ip4(
        n12900), .op(n12905) );
  nand2_1 U15774 ( .ip1(n13166), .ip2(n12903), .op(n12904) );
  nand3_1 U15775 ( .ip1(n12906), .ip2(n12905), .ip3(n12904), .op(n12907) );
  mux2_1 U15776 ( .ip1(data_wr_mem[16]), .ip2(n12907), .s(n13033), .op(n5272)
         );
  nand2_1 U15777 ( .ip1(n13172), .ip2(n12908), .op(n12924) );
  nor2_1 U15778 ( .ip1(n12909), .ip2(n13163), .op(n12919) );
  nand2_1 U15779 ( .ip1(n13162), .ip2(n12910), .op(n12917) );
  nand2_1 U15780 ( .ip1(n13180), .ip2(n12911), .op(n12916) );
  nand2_1 U15781 ( .ip1(n13168), .ip2(n12912), .op(n12915) );
  nand2_1 U15782 ( .ip1(n13170), .ip2(n12913), .op(n12914) );
  nand4_1 U15783 ( .ip1(n12917), .ip2(n12916), .ip3(n12915), .ip4(n12914), 
        .op(n12918) );
  not_ab_or_c_or_d U15784 ( .ip1(n13182), .ip2(n12920), .ip3(n12919), .ip4(
        n12918), .op(n12923) );
  nand2_1 U15785 ( .ip1(n13166), .ip2(n12921), .op(n12922) );
  nand3_1 U15786 ( .ip1(n12924), .ip2(n12923), .ip3(n12922), .op(n12925) );
  mux2_1 U15787 ( .ip1(data_wr_mem[17]), .ip2(n12925), .s(n13033), .op(n5271)
         );
  nand2_1 U15788 ( .ip1(n13170), .ip2(n12926), .op(n12942) );
  nor2_1 U15789 ( .ip1(n12927), .ip2(n13163), .op(n12937) );
  nand2_1 U15790 ( .ip1(n13168), .ip2(n12928), .op(n12935) );
  nand2_1 U15791 ( .ip1(n13182), .ip2(n12929), .op(n12934) );
  nand2_1 U15792 ( .ip1(n13172), .ip2(n12930), .op(n12933) );
  nand2_1 U15793 ( .ip1(n13162), .ip2(n12931), .op(n12932) );
  nand4_1 U15794 ( .ip1(n12935), .ip2(n12934), .ip3(n12933), .ip4(n12932), 
        .op(n12936) );
  not_ab_or_c_or_d U15795 ( .ip1(n13180), .ip2(n12938), .ip3(n12937), .ip4(
        n12936), .op(n12941) );
  nand2_1 U15796 ( .ip1(n13166), .ip2(n12939), .op(n12940) );
  nand3_1 U15797 ( .ip1(n12942), .ip2(n12941), .ip3(n12940), .op(n12943) );
  mux2_1 U15798 ( .ip1(data_wr_mem[18]), .ip2(n12943), .s(n13033), .op(n5270)
         );
  nand2_1 U15799 ( .ip1(n13168), .ip2(n12944), .op(n12960) );
  nor2_1 U15800 ( .ip1(n12945), .ip2(n13163), .op(n12955) );
  nand2_1 U15801 ( .ip1(n13170), .ip2(n12946), .op(n12953) );
  nand2_1 U15802 ( .ip1(n13172), .ip2(n12947), .op(n12952) );
  nand2_1 U15803 ( .ip1(n13182), .ip2(n12948), .op(n12951) );
  nand2_1 U15804 ( .ip1(n13180), .ip2(n12949), .op(n12950) );
  nand4_1 U15805 ( .ip1(n12953), .ip2(n12952), .ip3(n12951), .ip4(n12950), 
        .op(n12954) );
  not_ab_or_c_or_d U15806 ( .ip1(n13166), .ip2(n12956), .ip3(n12955), .ip4(
        n12954), .op(n12959) );
  nand2_1 U15807 ( .ip1(n13162), .ip2(n12957), .op(n12958) );
  nand3_1 U15808 ( .ip1(n12960), .ip2(n12959), .ip3(n12958), .op(n12961) );
  mux2_1 U15809 ( .ip1(data_wr_mem[19]), .ip2(n12961), .s(n13033), .op(n5269)
         );
  nand2_1 U15810 ( .ip1(n13180), .ip2(n12962), .op(n12978) );
  nor2_1 U15811 ( .ip1(n12963), .ip2(n13163), .op(n12973) );
  nand2_1 U15812 ( .ip1(n13182), .ip2(n12964), .op(n12971) );
  nand2_1 U15813 ( .ip1(n13162), .ip2(n12965), .op(n12970) );
  nand2_1 U15814 ( .ip1(n13172), .ip2(n12966), .op(n12969) );
  nand2_1 U15815 ( .ip1(n13170), .ip2(n12967), .op(n12968) );
  nand4_1 U15816 ( .ip1(n12971), .ip2(n12970), .ip3(n12969), .ip4(n12968), 
        .op(n12972) );
  not_ab_or_c_or_d U15817 ( .ip1(n13166), .ip2(n12974), .ip3(n12973), .ip4(
        n12972), .op(n12977) );
  nand2_1 U15818 ( .ip1(n13168), .ip2(n12975), .op(n12976) );
  nand3_1 U15819 ( .ip1(n12978), .ip2(n12977), .ip3(n12976), .op(n12979) );
  mux2_1 U15820 ( .ip1(data_wr_mem[20]), .ip2(n12979), .s(n13033), .op(n5268)
         );
  nand2_1 U15821 ( .ip1(n13170), .ip2(n12980), .op(n12996) );
  nor2_1 U15822 ( .ip1(n12981), .ip2(n13163), .op(n12991) );
  nand2_1 U15823 ( .ip1(n13180), .ip2(n12982), .op(n12989) );
  nand2_1 U15824 ( .ip1(n13172), .ip2(n12983), .op(n12988) );
  nand2_1 U15825 ( .ip1(n13168), .ip2(n12984), .op(n12987) );
  nand2_1 U15826 ( .ip1(n13166), .ip2(n12985), .op(n12986) );
  nand4_1 U15827 ( .ip1(n12989), .ip2(n12988), .ip3(n12987), .ip4(n12986), 
        .op(n12990) );
  not_ab_or_c_or_d U15828 ( .ip1(n13162), .ip2(n12992), .ip3(n12991), .ip4(
        n12990), .op(n12995) );
  nand2_1 U15829 ( .ip1(n13182), .ip2(n12993), .op(n12994) );
  nand3_1 U15830 ( .ip1(n12996), .ip2(n12995), .ip3(n12994), .op(n12997) );
  mux2_1 U15831 ( .ip1(data_wr_mem[21]), .ip2(n12997), .s(n13033), .op(n5267)
         );
  nand2_1 U15832 ( .ip1(n13168), .ip2(n12998), .op(n13014) );
  nor2_1 U15833 ( .ip1(n12999), .ip2(n13163), .op(n13009) );
  nand2_1 U15834 ( .ip1(n13172), .ip2(n13000), .op(n13007) );
  nand2_1 U15835 ( .ip1(n13180), .ip2(n13001), .op(n13006) );
  nand2_1 U15836 ( .ip1(n13166), .ip2(n13002), .op(n13005) );
  nand2_1 U15837 ( .ip1(n13170), .ip2(n13003), .op(n13004) );
  nand4_1 U15838 ( .ip1(n13007), .ip2(n13006), .ip3(n13005), .ip4(n13004), 
        .op(n13008) );
  not_ab_or_c_or_d U15839 ( .ip1(n13182), .ip2(n13010), .ip3(n13009), .ip4(
        n13008), .op(n13013) );
  nand2_1 U15840 ( .ip1(n13162), .ip2(n13011), .op(n13012) );
  nand3_1 U15841 ( .ip1(n13014), .ip2(n13013), .ip3(n13012), .op(n13015) );
  mux2_1 U15842 ( .ip1(data_wr_mem[22]), .ip2(n13015), .s(n13033), .op(n5266)
         );
  nand2_1 U15843 ( .ip1(n13172), .ip2(n13016), .op(n13032) );
  nor2_1 U15844 ( .ip1(n13017), .ip2(n13163), .op(n13027) );
  nand2_1 U15845 ( .ip1(n13162), .ip2(n13018), .op(n13025) );
  nand2_1 U15846 ( .ip1(n13180), .ip2(n13019), .op(n13024) );
  nand2_1 U15847 ( .ip1(n13182), .ip2(n13020), .op(n13023) );
  nand2_1 U15848 ( .ip1(n13166), .ip2(n13021), .op(n13022) );
  nand4_1 U15849 ( .ip1(n13025), .ip2(n13024), .ip3(n13023), .ip4(n13022), 
        .op(n13026) );
  not_ab_or_c_or_d U15850 ( .ip1(n13170), .ip2(n13028), .ip3(n13027), .ip4(
        n13026), .op(n13031) );
  nand2_1 U15851 ( .ip1(n13168), .ip2(n13029), .op(n13030) );
  nand3_1 U15852 ( .ip1(n13032), .ip2(n13031), .ip3(n13030), .op(n13034) );
  mux2_1 U15853 ( .ip1(data_wr_mem[23]), .ip2(n13034), .s(n13033), .op(n5265)
         );
  nand2_1 U15854 ( .ip1(n13180), .ip2(n13035), .op(n13051) );
  nor2_1 U15855 ( .ip1(n13036), .ip2(n13163), .op(n13046) );
  nand2_1 U15856 ( .ip1(n13166), .ip2(n13037), .op(n13044) );
  nand2_1 U15857 ( .ip1(n13170), .ip2(n13038), .op(n13043) );
  nand2_1 U15858 ( .ip1(n13182), .ip2(n13039), .op(n13042) );
  nand2_1 U15859 ( .ip1(n13172), .ip2(n13040), .op(n13041) );
  nand4_1 U15860 ( .ip1(n13044), .ip2(n13043), .ip3(n13042), .ip4(n13041), 
        .op(n13045) );
  not_ab_or_c_or_d U15861 ( .ip1(n13162), .ip2(n13047), .ip3(n13046), .ip4(
        n13045), .op(n13050) );
  nand2_1 U15862 ( .ip1(n13168), .ip2(n13048), .op(n13049) );
  nand3_1 U15863 ( .ip1(n13051), .ip2(n13050), .ip3(n13049), .op(n13052) );
  mux2_1 U15864 ( .ip1(data_wr_mem[24]), .ip2(n13052), .s(n13186), .op(n5264)
         );
  nand2_1 U15865 ( .ip1(n13182), .ip2(n13053), .op(n13069) );
  nor2_1 U15866 ( .ip1(n13054), .ip2(n13163), .op(n13064) );
  nand2_1 U15867 ( .ip1(n13170), .ip2(n13055), .op(n13062) );
  nand2_1 U15868 ( .ip1(n13180), .ip2(n13056), .op(n13061) );
  nand2_1 U15869 ( .ip1(n13162), .ip2(n13057), .op(n13060) );
  nand2_1 U15870 ( .ip1(n13168), .ip2(n13058), .op(n13059) );
  nand4_1 U15871 ( .ip1(n13062), .ip2(n13061), .ip3(n13060), .ip4(n13059), 
        .op(n13063) );
  not_ab_or_c_or_d U15872 ( .ip1(n13172), .ip2(n13065), .ip3(n13064), .ip4(
        n13063), .op(n13068) );
  nand2_1 U15873 ( .ip1(n13166), .ip2(n13066), .op(n13067) );
  nand3_1 U15874 ( .ip1(n13069), .ip2(n13068), .ip3(n13067), .op(n13070) );
  mux2_1 U15875 ( .ip1(data_wr_mem[25]), .ip2(n13070), .s(n13186), .op(n5263)
         );
  nand2_1 U15876 ( .ip1(n13168), .ip2(n13071), .op(n13087) );
  nor2_1 U15877 ( .ip1(n13072), .ip2(n13163), .op(n13082) );
  nand2_1 U15878 ( .ip1(n13162), .ip2(n13073), .op(n13080) );
  nand2_1 U15879 ( .ip1(n13172), .ip2(n13074), .op(n13079) );
  nand2_1 U15880 ( .ip1(n13180), .ip2(n13075), .op(n13078) );
  nand2_1 U15881 ( .ip1(n13166), .ip2(n13076), .op(n13077) );
  nand4_1 U15882 ( .ip1(n13080), .ip2(n13079), .ip3(n13078), .ip4(n13077), 
        .op(n13081) );
  not_ab_or_c_or_d U15883 ( .ip1(n13170), .ip2(n13083), .ip3(n13082), .ip4(
        n13081), .op(n13086) );
  nand2_1 U15884 ( .ip1(n13182), .ip2(n13084), .op(n13085) );
  nand3_1 U15885 ( .ip1(n13087), .ip2(n13086), .ip3(n13085), .op(n13088) );
  mux2_1 U15886 ( .ip1(data_wr_mem[26]), .ip2(n13088), .s(n13186), .op(n5262)
         );
  nand2_1 U15887 ( .ip1(n13168), .ip2(n13089), .op(n13105) );
  nor2_1 U15888 ( .ip1(n13090), .ip2(n13163), .op(n13100) );
  nand2_1 U15889 ( .ip1(n13166), .ip2(n13091), .op(n13098) );
  nand2_1 U15890 ( .ip1(n13172), .ip2(n13092), .op(n13097) );
  nand2_1 U15891 ( .ip1(n13180), .ip2(n13093), .op(n13096) );
  nand2_1 U15892 ( .ip1(n13170), .ip2(n13094), .op(n13095) );
  nand4_1 U15893 ( .ip1(n13098), .ip2(n13097), .ip3(n13096), .ip4(n13095), 
        .op(n13099) );
  not_ab_or_c_or_d U15894 ( .ip1(n13182), .ip2(n13101), .ip3(n13100), .ip4(
        n13099), .op(n13104) );
  nand2_1 U15895 ( .ip1(n13162), .ip2(n13102), .op(n13103) );
  nand3_1 U15896 ( .ip1(n13105), .ip2(n13104), .ip3(n13103), .op(n13106) );
  mux2_1 U15897 ( .ip1(data_wr_mem[27]), .ip2(n13106), .s(n13186), .op(n5261)
         );
  nand2_1 U15898 ( .ip1(n13168), .ip2(n13107), .op(n13123) );
  nor2_1 U15899 ( .ip1(n13108), .ip2(n13163), .op(n13118) );
  nand2_1 U15900 ( .ip1(n13166), .ip2(n13109), .op(n13116) );
  nand2_1 U15901 ( .ip1(n13172), .ip2(n13110), .op(n13115) );
  nand2_1 U15902 ( .ip1(n13180), .ip2(n13111), .op(n13114) );
  nand2_1 U15903 ( .ip1(n13170), .ip2(n13112), .op(n13113) );
  nand4_1 U15904 ( .ip1(n13116), .ip2(n13115), .ip3(n13114), .ip4(n13113), 
        .op(n13117) );
  not_ab_or_c_or_d U15905 ( .ip1(n13162), .ip2(n13119), .ip3(n13118), .ip4(
        n13117), .op(n13122) );
  nand2_1 U15906 ( .ip1(n13182), .ip2(n13120), .op(n13121) );
  nand3_1 U15907 ( .ip1(n13123), .ip2(n13122), .ip3(n13121), .op(n13124) );
  mux2_1 U15908 ( .ip1(data_wr_mem[28]), .ip2(n13124), .s(n13186), .op(n5260)
         );
  nand2_1 U15909 ( .ip1(n13166), .ip2(n13125), .op(n13141) );
  nor2_1 U15910 ( .ip1(n13126), .ip2(n13163), .op(n13136) );
  nand2_1 U15911 ( .ip1(n13170), .ip2(n13127), .op(n13134) );
  nand2_1 U15912 ( .ip1(n13180), .ip2(n13128), .op(n13133) );
  nand2_1 U15913 ( .ip1(n13168), .ip2(n13129), .op(n13132) );
  nand2_1 U15914 ( .ip1(n13172), .ip2(n13130), .op(n13131) );
  nand4_1 U15915 ( .ip1(n13134), .ip2(n13133), .ip3(n13132), .ip4(n13131), 
        .op(n13135) );
  not_ab_or_c_or_d U15916 ( .ip1(n13182), .ip2(n13137), .ip3(n13136), .ip4(
        n13135), .op(n13140) );
  nand2_1 U15917 ( .ip1(n13162), .ip2(n13138), .op(n13139) );
  nand3_1 U15918 ( .ip1(n13141), .ip2(n13140), .ip3(n13139), .op(n13142) );
  mux2_1 U15919 ( .ip1(data_wr_mem[29]), .ip2(n13142), .s(n13186), .op(n5259)
         );
  nand2_1 U15920 ( .ip1(n13162), .ip2(n13143), .op(n13159) );
  nor2_1 U15921 ( .ip1(n13144), .ip2(n13163), .op(n13154) );
  nand2_1 U15922 ( .ip1(n13166), .ip2(n13145), .op(n13152) );
  nand2_1 U15923 ( .ip1(n13180), .ip2(n13146), .op(n13151) );
  nand2_1 U15924 ( .ip1(n13168), .ip2(n13147), .op(n13150) );
  nand2_1 U15925 ( .ip1(n13170), .ip2(n13148), .op(n13149) );
  nand4_1 U15926 ( .ip1(n13152), .ip2(n13151), .ip3(n13150), .ip4(n13149), 
        .op(n13153) );
  not_ab_or_c_or_d U15927 ( .ip1(n13172), .ip2(n13155), .ip3(n13154), .ip4(
        n13153), .op(n13158) );
  nand2_1 U15928 ( .ip1(n13182), .ip2(n13156), .op(n13157) );
  nand3_1 U15929 ( .ip1(n13159), .ip2(n13158), .ip3(n13157), .op(n13160) );
  mux2_1 U15930 ( .ip1(data_wr_mem[30]), .ip2(n13160), .s(n13186), .op(n5258)
         );
  nand2_1 U15931 ( .ip1(n13162), .ip2(n13161), .op(n13185) );
  nor2_1 U15932 ( .ip1(n13164), .ip2(n13163), .op(n13178) );
  nand2_1 U15933 ( .ip1(n13166), .ip2(n13165), .op(n13176) );
  nand2_1 U15934 ( .ip1(n13168), .ip2(n13167), .op(n13175) );
  nand2_1 U15935 ( .ip1(n13170), .ip2(n13169), .op(n13174) );
  nand2_1 U15936 ( .ip1(n13172), .ip2(n13171), .op(n13173) );
  nand4_1 U15937 ( .ip1(n13176), .ip2(n13175), .ip3(n13174), .ip4(n13173), 
        .op(n13177) );
  not_ab_or_c_or_d U15938 ( .ip1(n13180), .ip2(n13179), .ip3(n13178), .ip4(
        n13177), .op(n13184) );
  nand2_1 U15939 ( .ip1(n13182), .ip2(n13181), .op(n13183) );
  nand3_1 U15940 ( .ip1(n13185), .ip2(n13184), .ip3(n13183), .op(n13187) );
  mux2_1 U15941 ( .ip1(data_wr_mem[31]), .ip2(n13187), .s(n13186), .op(n5257)
         );
  nand2_1 U15942 ( .ip1(wr_mem), .ip2(n13201), .op(n13188) );
  nand2_1 U15943 ( .ip1(n13189), .ip2(n13188), .op(n5256) );
  nand2_1 U15944 ( .ip1(rd_mem), .ip2(n13201), .op(n13190) );
  nand2_1 U15945 ( .ip1(n13191), .ip2(n13190), .op(n5255) );
  nand2_1 U15946 ( .ip1(addr_mem[2]), .ip2(n13201), .op(n13192) );
  nand2_1 U15947 ( .ip1(n13193), .ip2(n13192), .op(n5252) );
  nand2_1 U15948 ( .ip1(mem_data_cnt[3]), .ip2(n13200), .op(n13195) );
  nand2_1 U15949 ( .ip1(addr_mem[3]), .ip2(n13201), .op(n13194) );
  nand2_1 U15950 ( .ip1(n13195), .ip2(n13194), .op(n5251) );
  nand2_1 U15951 ( .ip1(addr_resp[4]), .ip2(n13200), .op(n13197) );
  nand2_1 U15952 ( .ip1(addr_mem[4]), .ip2(n13201), .op(n13196) );
  nand2_1 U15953 ( .ip1(n13197), .ip2(n13196), .op(n5250) );
  nand2_1 U15954 ( .ip1(addr_resp[5]), .ip2(n13200), .op(n13199) );
  nand2_1 U15955 ( .ip1(addr_mem[5]), .ip2(n13201), .op(n13198) );
  nand2_1 U15956 ( .ip1(n13199), .ip2(n13198), .op(n5249) );
  nand2_1 U15957 ( .ip1(addr_resp[6]), .ip2(n13200), .op(n13203) );
  nand2_1 U15958 ( .ip1(addr_mem[6]), .ip2(n13201), .op(n13202) );
  nand2_1 U15959 ( .ip1(n13203), .ip2(n13202), .op(n5248) );
  nand2_1 U15961 ( .ip1(miss), .ip2(n13290), .op(n13204) );
  nand2_1 U15962 ( .ip1(n13205), .ip2(n13204), .op(n5221) );
  nand2_1 U15963 ( .ip1(n13209), .ip2(cache_miss_count[29]), .op(n13207) );
  inv_1 U15964 ( .ip(cache_miss_count[30]), .op(n13208) );
  nor2_1 U15965 ( .ip1(n13207), .ip2(n13208), .op(n13206) );
  xor2_1 U15966 ( .ip1(n13206), .ip2(cache_miss_count[31]), .op(n5220) );
  mux2_1 U15967 ( .ip1(n13208), .ip2(cache_miss_count[30]), .s(n13207), .op(
        n5219) );
  xor2_1 U15968 ( .ip1(n13209), .ip2(cache_miss_count[29]), .op(n5218) );
  xor2_1 U15969 ( .ip1(n13210), .ip2(cache_miss_count[27]), .op(n5216) );
  xor2_1 U15970 ( .ip1(n13211), .ip2(cache_miss_count[25]), .op(n5214) );
  xor2_1 U15971 ( .ip1(n13212), .ip2(cache_miss_count[23]), .op(n5212) );
  xor2_1 U15972 ( .ip1(n13213), .ip2(cache_miss_count[21]), .op(n5210) );
  xor2_1 U15973 ( .ip1(n13214), .ip2(cache_miss_count[19]), .op(n5208) );
  xor2_1 U15974 ( .ip1(n13215), .ip2(cache_miss_count[17]), .op(n5206) );
  xor2_1 U15975 ( .ip1(n13216), .ip2(cache_miss_count[15]), .op(n5204) );
  xor2_1 U15976 ( .ip1(n13217), .ip2(cache_miss_count[13]), .op(n5202) );
  xor2_1 U15977 ( .ip1(n13218), .ip2(cache_miss_count[11]), .op(n5200) );
  inv_1 U15978 ( .ip(cache_miss_count[9]), .op(n13220) );
  mux2_1 U15979 ( .ip1(cache_miss_count[9]), .ip2(n13220), .s(n13219), .op(
        n5198) );
  mux2_1 U15980 ( .ip1(n13224), .ip2(n13221), .s(cache_miss_count[7]), .op(
        n5196) );
  nor2_1 U15981 ( .ip1(n13222), .ip2(cache_miss_count[6]), .op(n13223) );
  nor2_1 U15982 ( .ip1(n13224), .ip2(n13223), .op(n5195) );
  inv_1 U15983 ( .ip(cache_miss_count[4]), .op(n13226) );
  mux2_1 U15984 ( .ip1(cache_miss_count[4]), .ip2(n13226), .s(n13225), .op(
        n5193) );
  inv_1 U15985 ( .ip(n13227), .op(n13230) );
  nor2_1 U15986 ( .ip1(n13228), .ip2(cache_miss_count[2]), .op(n13229) );
  nor2_1 U15987 ( .ip1(n13230), .ip2(n13229), .op(n5191) );
  inv_1 U15988 ( .ip(n13231), .op(n13232) );
  mux2_1 U15989 ( .ip1(n13232), .ip2(n13231), .s(cache_miss_count[0]), .op(
        n5189) );
  nand2_1 U15990 ( .ip1(n13236), .ip2(cache_hit_count[29]), .op(n13234) );
  inv_1 U15991 ( .ip(cache_hit_count[30]), .op(n13235) );
  nor2_1 U15992 ( .ip1(n13234), .ip2(n13235), .op(n13233) );
  xor2_1 U15993 ( .ip1(n13233), .ip2(cache_hit_count[31]), .op(n5187) );
  mux2_1 U15994 ( .ip1(n13235), .ip2(cache_hit_count[30]), .s(n13234), .op(
        n5186) );
  xor2_1 U15995 ( .ip1(n13236), .ip2(cache_hit_count[29]), .op(n5185) );
  xor2_1 U15996 ( .ip1(n13237), .ip2(cache_hit_count[27]), .op(n5183) );
  xor2_1 U15997 ( .ip1(n13238), .ip2(cache_hit_count[25]), .op(n5181) );
  xor2_1 U15998 ( .ip1(n13239), .ip2(cache_hit_count[23]), .op(n5179) );
  xor2_1 U15999 ( .ip1(n13240), .ip2(cache_hit_count[21]), .op(n5177) );
  xor2_1 U16000 ( .ip1(n13241), .ip2(cache_hit_count[19]), .op(n5175) );
  xor2_1 U16001 ( .ip1(n13242), .ip2(cache_hit_count[17]), .op(n5173) );
  xor2_1 U16002 ( .ip1(n13243), .ip2(cache_hit_count[15]), .op(n5171) );
  xor2_1 U16003 ( .ip1(n13244), .ip2(cache_hit_count[13]), .op(n5169) );
  xor2_1 U16004 ( .ip1(n13245), .ip2(cache_hit_count[11]), .op(n5167) );
  xor2_1 U16005 ( .ip1(n13246), .ip2(cache_hit_count[9]), .op(n5165) );
  xor2_1 U16006 ( .ip1(n13247), .ip2(cache_hit_count[7]), .op(n5163) );
  xor2_1 U16007 ( .ip1(n13248), .ip2(cache_hit_count[5]), .op(n5161) );
  xor2_1 U16008 ( .ip1(n13249), .ip2(cache_hit_count[3]), .op(n5159) );
  xor2_1 U16009 ( .ip1(n13250), .ip2(cache_hit_count[1]), .op(n5157) );
  nand2_1 U16010 ( .ip1(n13251), .ip2(cache_valid_A[6]), .op(n13263) );
  nor2_1 U16011 ( .ip1(n9178), .ip2(n13252), .op(n13260) );
  nand2_1 U16012 ( .ip1(n13253), .ip2(cache_valid_A[3]), .op(n13258) );
  nand2_1 U16013 ( .ip1(n13254), .ip2(cache_valid_A[5]), .op(n13257) );
  nand2_1 U16014 ( .ip1(n13270), .ip2(cache_valid_A[0]), .op(n13256) );
  nand2_1 U16015 ( .ip1(n13278), .ip2(cache_valid_A[1]), .op(n13255) );
  nand4_1 U16016 ( .ip1(n13258), .ip2(n13257), .ip3(n13256), .ip4(n13255), 
        .op(n13259) );
  not_ab_or_c_or_d U16017 ( .ip1(n13264), .ip2(cache_valid_A[2]), .ip3(n13260), 
        .ip4(n13259), .op(n13262) );
  nand2_1 U16018 ( .ip1(n13268), .ip2(cache_valid_A[4]), .op(n13261) );
  nand3_1 U16019 ( .ip1(n13263), .ip2(n13262), .ip3(n13261), .op(n13289) );
  nand2_1 U16020 ( .ip1(cache_valid_B[2]), .ip2(n13264), .op(n13281) );
  nor2_1 U16021 ( .ip1(n13266), .ip2(n13265), .op(n13276) );
  nand2_1 U16022 ( .ip1(n13267), .ip2(cache_valid_B[5]), .op(n13274) );
  nand2_1 U16023 ( .ip1(n13268), .ip2(cache_valid_B[4]), .op(n13273) );
  nand2_1 U16024 ( .ip1(n13269), .ip2(cache_valid_B[6]), .op(n13272) );
  nand2_1 U16025 ( .ip1(n13270), .ip2(cache_valid_B[0]), .op(n13271) );
  nand4_1 U16026 ( .ip1(n13274), .ip2(n13273), .ip3(n13272), .ip4(n13271), 
        .op(n13275) );
  not_ab_or_c_or_d U16027 ( .ip1(cache_valid_B[7]), .ip2(n13277), .ip3(n13276), 
        .ip4(n13275), .op(n13280) );
  nand2_1 U16028 ( .ip1(n13278), .ip2(cache_valid_B[1]), .op(n13279) );
  nand3_1 U16029 ( .ip1(n13281), .ip2(n13280), .ip3(n13279), .op(n13288) );
  or2_1 U16030 ( .ip1(n13282), .ip2(n13283), .op(n13286) );
  or2_1 U16031 ( .ip1(n13284), .ip2(n13283), .op(n13285) );
  nand2_1 U16032 ( .ip1(n13286), .ip2(n13285), .op(n13287) );
  mux2_1 U16033 ( .ip1(n13289), .ip2(n13288), .s(n13287), .op(n13291) );
  mux2_1 U16034 ( .ip1(n13291), .ip2(valid), .s(n13290), .op(n5155) );
  inv_1 U16035 ( .ip(N4300), .op(n127) );
  inv_1 U16036 ( .ip(N4297), .op(n125) );
  inv_1 U16037 ( .ip(N4294), .op(n123) );
  inv_1 U16038 ( .ip(N4291), .op(n121) );
  inv_1 U16039 ( .ip(N4288), .op(n119) );
  inv_1 U16040 ( .ip(N4285), .op(n117) );
  inv_1 U16041 ( .ip(N4282), .op(n115) );
  inv_1 U16042 ( .ip(N4279), .op(n113) );
  inv_1 U16043 ( .ip(N4276), .op(n111) );
  inv_1 U16044 ( .ip(N4273), .op(n109) );
  inv_1 U16045 ( .ip(N4270), .op(n107) );
  inv_1 U16046 ( .ip(N4267), .op(n105) );
  inv_1 U16047 ( .ip(N4264), .op(n103) );
  inv_1 U16048 ( .ip(N4261), .op(n101) );
  inv_1 U16049 ( .ip(N4258), .op(n99) );
  inv_1 U16050 ( .ip(N4255), .op(n97) );
  inv_1 U16051 ( .ip(N4252), .op(n95) );
  inv_1 U16052 ( .ip(N4249), .op(n93) );
  inv_1 U16053 ( .ip(N4246), .op(n91) );
  inv_1 U16054 ( .ip(N4243), .op(n89) );
  inv_1 U16055 ( .ip(N4240), .op(n87) );
  inv_1 U16056 ( .ip(N4237), .op(n85) );
  inv_1 U16057 ( .ip(N4234), .op(n83) );
  inv_1 U16058 ( .ip(N4231), .op(n81) );
  inv_1 U16059 ( .ip(N4228), .op(n79) );
  inv_1 U16060 ( .ip(N4225), .op(n77) );
  inv_1 U16061 ( .ip(N4222), .op(n75) );
  inv_1 U16062 ( .ip(N4219), .op(n73) );
  inv_1 U16063 ( .ip(N4216), .op(n71) );
  inv_1 U16064 ( .ip(N4213), .op(n69) );
  inv_1 U16065 ( .ip(N4210), .op(n67) );
  inv_1 U16066 ( .ip(N4207), .op(n65) );
  inv_1 U16067 ( .ip(N4204), .op(n63) );
  inv_1 U16068 ( .ip(N4201), .op(n61) );
  inv_1 U16069 ( .ip(N4198), .op(n59) );
  inv_1 U16070 ( .ip(N4195), .op(n57) );
  inv_1 U16071 ( .ip(N4192), .op(n55) );
  inv_1 U16072 ( .ip(N4189), .op(n53) );
  inv_1 U16073 ( .ip(N4186), .op(n51) );
  inv_1 U16074 ( .ip(N4183), .op(n49) );
  inv_1 U16075 ( .ip(N4180), .op(n47) );
  inv_1 U16076 ( .ip(N4177), .op(n45) );
  inv_1 U16077 ( .ip(N4174), .op(n43) );
  inv_1 U16078 ( .ip(N4171), .op(n41) );
  inv_1 U16079 ( .ip(N4168), .op(n39) );
  inv_1 U16080 ( .ip(N4165), .op(n37) );
  inv_1 U16081 ( .ip(N4162), .op(n35) );
  inv_1 U16082 ( .ip(N4159), .op(n33) );
  inv_1 U16083 ( .ip(N4156), .op(n31) );
  inv_1 U16084 ( .ip(N4153), .op(n29) );
  inv_1 U16085 ( .ip(N4150), .op(n27) );
  inv_1 U16086 ( .ip(N4147), .op(n25) );
  inv_1 U16087 ( .ip(N4144), .op(n23) );
  inv_1 U16088 ( .ip(N4141), .op(n21) );
  inv_1 U16089 ( .ip(N4138), .op(n19) );
  inv_1 U16090 ( .ip(N4135), .op(n17) );
  inv_1 U16091 ( .ip(N4132), .op(n15) );
  inv_1 U16092 ( .ip(N4129), .op(n13) );
  inv_1 U16093 ( .ip(N4126), .op(n11) );
  inv_1 U16094 ( .ip(N4123), .op(n9) );
  inv_1 U16095 ( .ip(N4120), .op(n7) );
  inv_1 U16096 ( .ip(N4117), .op(n5) );
  inv_1 U16097 ( .ip(N4114), .op(n3) );
  inv_1 U16098 ( .ip(N4111), .op(n1) );
endmodule

